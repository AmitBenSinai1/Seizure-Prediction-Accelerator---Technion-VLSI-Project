/*------------------------------------------------------------------------------
 * File          : define.sv
 * Project       : RTL
 * Author        : epamof
 * Creation date : Mar 10, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

`define FIFO_ADDR 10'h0
`define FIFO_DATA 10'h1
`define START_ADDR 10'h2

`define LUT_ADDR 10'h3
`define LUT_DATA_1 10'h4
`define LUT_DATA_2 10'h5
`define LUT_DATA_3 10'h6


`define NUM_OF_INPUTS 9'100000000 // 256

