/*------------------------------------------------------------------------------
 * File          : seizure_tb.sv
 * Project       : RTL
 * Author        : epamof
 * Creation date : Feb 15, 2024
 * Description   :
 *------------------------------------------------------------------------------*/
`timescale 1ns/1ps
`include "/users/epamof/Project/design/define.sv"
//`include "/users/epamof/Project/design/write_lut_mcmc.sv"

module seizure_tb #() ();

// Constants
parameter CLK_PERIOD = 10; // Clock period in nanoseconds

// Signals
logic apb_clk;
logic reset_n;
logic [9:0] apb_addr = `FIFO_DATA;
logic apb_psel;
logic apb_penable;
logic apb_pwrite;
logic [31:0] apb_pwdata;
logic [31:0] apb_prdata;
logic apb_ready;
logic [31:0] read_reg_data;
logic [17:0] read_fifo_data;
logic seizure_prediction;


// Instantiate the seizure_top module
seizure_top seizure_top (
	.apb_clk(apb_clk),
	.reset_n(reset_n),
	.apb_addr(apb_addr),
	.apb_pwrite(apb_pwrite),
	.apb_psel(apb_psel),
	.apb_penable(apb_penable),
	.apb_pwdata(apb_pwdata),
	.apb_prdata(apb_prdata),
	.apb_ready(apb_ready),
	.seizure_prediction(seizure_prediction)
);

// Clock generation
always begin
	#(CLK_PERIOD/2) apb_clk = ~apb_clk;
end

// Task to perform APB write
task apb_write(input logic [9:0] addr, input logic [31:0] data);
	begin
		apb_addr = addr;
		apb_penable = 1;
		apb_pwrite = 1; // Write operation
		apb_pwdata = data; // Write data
		#10 apb_penable = 0; // Deassert peripheral enable
	end
endtask

// Task to perform APB read
task apb_read(input logic [9:0] addr);
	begin
		apb_addr = addr;
		apb_penable = 1;
		apb_pwrite = 0; // Read operation
		#10 apb_penable = 0; // Deassert peripheral enable
		read_reg_data = apb_prdata; // Capture read data
		$display("APB read: address=%s, data=%s", addr, read_reg_data);
	end
endtask



task FIFO_indirect_write(input logic [7:0] addr,  input logic [17:0] data);
	begin
		apb_write(`FIFO_ADDR, addr);
		apb_write(`FIFO_DATA, data);
	end
endtask
	
	
task FIFO_indirect_read(input logic [7:0] addr);
	begin
		apb_write(`FIFO_ADDR, addr);
		apb_read(`FIFO_DATA);
	end
endtask

///////////////////



task MCMC_indirect_write(input logic [10:0] addr,  input logic [67:0] data);
	begin
		apb_write(`LUT_ADDR, addr);
		apb_write(`LUT_DATA_1, data[67:64]);
		apb_write(`LUT_DATA_2, data[63:32]);
		apb_write(`LUT_DATA_3, data[31:0]);
	end
endtask
	
	
task MCMC_indirect_read(input logic [10:0] addr);
	begin
		apb_write(`LUT_ADDR, addr);
		apb_read(`LUT_DATA_3);
		apb_read(`LUT_DATA_2);
		apb_read(`LUT_DATA_1);
	end
endtask
///////////////
// Test stimulus
initial begin
	apb_clk = 0;
	reset_n = 0; // Assert reset
	apb_addr = 10'b0;
	apb_pwrite = 0;
	apb_psel = 1;
	apb_pwdata = 32'h0;
	apb_penable = 1'b0;
	#100 reset_n = 1; // Deassert reset after 100 time units

	//pc
	//indirect write - 256 times
	//start_pc - start count
	
	FIFO_indirect_write(8'd0, 18'b000000100000000000); #20	// 1  EEG signal     0 00000 1000 0000 0000 +0.5 || 800
	FIFO_indirect_write(8'd1, 18'b100010000000000000); #20	// 2  EEG signal     1 00010 0000 0000 0000 -2 || 2_2000
	FIFO_indirect_write(8'd2, 18'b000000010000000000); #20	// 3  EEG signal     0 00000 0100 0000 0000 +0.25 || 400
	FIFO_indirect_write(8'd3, 18'b101000100000000000); #20	// 4  EEG signal     1 01000 1000 0000 0000  -8.5 || 2_8800
			
	FIFO_indirect_write(8'd4, 18'b000000100000000000); #20	// 5  EEG signal     0 00000 1000 0000 0000 +0.5 || 800
	FIFO_indirect_write(8'd5, 18'b100010000000000000); #20	// 6  EEG signal     1 00010 0000 0000 0000 -2 || 2_2000
	FIFO_indirect_write(8'd6, 18'b000000010000000000); #20 	// 7  EEG signal     0 00000 0100 0000 0000 +0.25 || 400
	FIFO_indirect_write(8'd7, 18'b101000100000000000); #20 	// 8  EEG signal     1 01000 1000 0000 0000  -8.5 || 2_8800
							
	FIFO_indirect_write(8'd8, 18'b000011100000000000); #20	// 9  EEG signal   	 0 00011 1000 0000 0000 +3.5 || 3800
	FIFO_indirect_write(8'd9, 18'b100010110000000000); #20	// 10 EEG signal     1 00010 1100 0000 0000 -2.75 || 2_2c00
	FIFO_indirect_write(8'd10, 18'b010000010000000000); #20	// 11 EEG signal     0 10000 0100 0000 0000 +16.25 || 1_0400
	FIFO_indirect_write(8'd11, 18'b101000110000000000); #20	// 12 EEG signal     1 01000 1100 0000 0000  -8.75 || 2_8c00
			
	FIFO_indirect_write(8'd12, 18'b000000001000000000); #20	// 13 EEG signal     0 00000 0010 0000 0000 +0.125 || 200
	FIFO_indirect_write(8'd13, 18'b100010000000000000); #20	// 14 EEG signal     1 00010 0000 0000 0000 -2 || 2_2000
	FIFO_indirect_write(8'd14, 18'b000001010000000000); #20	// 15 EEG signal     0 00001 0100 0000 0000 +1.25 || 1400
	FIFO_indirect_write(8'd15, 18'b101000100000000000); #20	// 16 EEG signal     1 01000 1000 0000 0000  -8.5 || 2_8800
			
	
	// for dctc
	FIFO_indirect_write(8'd16, 18'b000001000000000000); #20	// 1  EEG signal     0 00001 0000 0000 0000 +1
	FIFO_indirect_write(8'd17, 18'b100001000000000000); #20	// 1  EEG signal     1 00001 0000 0000 0000 -1
	FIFO_indirect_write(8'd18, 18'b000010000000000000); #20	// 1  EEG signal     0 00010 0000 0000 0000 +2
	FIFO_indirect_write(8'd19, 18'b100010000000000000); #20	// 1  EEG signal     1 00010 0000 0000 0000 -2
	FIFO_indirect_write(8'd20, 18'b000011000000000000); #20	// 1  EEG signal     0 00011 0000 0000 0000 +3
	FIFO_indirect_write(8'd21, 18'b101000000000000000); #20	// 1  EEG signal     1 01000 0000 0000 0000 -8
	FIFO_indirect_write(8'd22, 18'b001100000000000000); #20	// 1  EEG signal     0 01100 0000 0000 0000 +12
	FIFO_indirect_write(8'd23, 18'b101000000000000000); #20	// 1  EEG signal     1 01000 0000 0000 0000 -8
	FIFO_indirect_write(8'd24, 18'b000000000000000000); #40	// 1  EEG signal     0 00000 0000 0000 0000 0
											


	
	/////////////////////
	
	MCMC_indirect_write(11'd0, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1, 68'b	00000010000110001000001010100001110000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd2, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd3, 68'b00000000000000000000000000000000000000000000000000000000101000110111); #20
	MCMC_indirect_write(11'd4, 68'b00101100001111111001010011010000010010110100000010100010111010001011); #20
	MCMC_indirect_write(11'd5, 68'b00100011010111010000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd6, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd7, 68'b00001011111000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd8, 68'b00010011011101100010000000010110110001011001000110000100111010001110); #20
	MCMC_indirect_write(11'd9, 68'b00101001110011010000111011010111000010000100001000000100001101111011); #20
	MCMC_indirect_write(11'd10, 68'b00000000000000000000100000101101110000111010100000100001100000011000); #20
	MCMC_indirect_write(11'd11, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd12, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd13, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd14, 68'b00000000000000000000000000000000000001110110100110100100010000011111); #20
	MCMC_indirect_write(11'd15, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd16, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd17, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd18, 68'b00100001010011001001000111010011010001000011111100100000000000000000); #20
	MCMC_indirect_write(11'd19, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd20, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd21, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd22, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd23, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd24, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd25, 68'b00000110011001101000010110001000110001001010011001100010001111110000); #20
	MCMC_indirect_write(11'd26, 68'b00101110100000011001010010100011100000010101000010100100110000111010); #20
	MCMC_indirect_write(11'd27, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd28, 68'b01010101101101110011001010111101000011110001111100001001101000010011); #20
	MCMC_indirect_write(11'd29, 68'b00001011110101101000000000000000000001111100111110000100000000100010); #20
	MCMC_indirect_write(11'd30, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd31, 68'b00011111000110111000011110001100100001101010110000100000000000000000); #20
	MCMC_indirect_write(11'd32, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd33, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd34, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd35, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd36, 68'b00000000000000000000000000000000000001110101100000100101001011110010); #20
	MCMC_indirect_write(11'd37, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd38, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd39, 68'b00000000000000000000000000000000000000001010110111100000000000000000); #20
	MCMC_indirect_write(11'd40, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd41, 68'b00000001010011110000000000000000000000101101000111100100110011101101); #20
	MCMC_indirect_write(11'd42, 68'b01000010010010111011010101111001010111010101001111001101111010110010); #20
	MCMC_indirect_write(11'd43, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd44, 68'b00001111100101011001010110101000010001010110011111100101100101110000); #20
	MCMC_indirect_write(11'd45, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd46, 68'b00000000000000000000000100001100010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd47, 68'b01100111111011101011100110100100110111100001011111010101011110100100); #20
	MCMC_indirect_write(11'd48, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd49, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd50, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd51, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd52, 68'b00101001101101101001101101101100100011000010011011000111101111000111); #20
	MCMC_indirect_write(11'd53, 68'b00111111011100000010100000010101110010101111010111100101101110001001); #20
	MCMC_indirect_write(11'd54, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd55, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd56, 68'b00000000000000000000011010011111010010101000001110100010111111011001); #20
	MCMC_indirect_write(11'd57, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd58, 68'b01000000110110011010010111010100000101011011111111001010110010110111); #20
	MCMC_indirect_write(11'd59, 68'b01100011110100110011101011010011100111111101110111001111111101101010); #20
	MCMC_indirect_write(11'd60, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd61, 68'b00000000000000000000000000000000000000111100101000100000001100101011); #20
	MCMC_indirect_write(11'd62, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd63, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd64, 68'b00001000000000000000010000000000000000100000000000000001000000000000); #20
	MCMC_indirect_write(11'd65, 68'b00000011101111110000001010100000100001001101010111100010000100100010); #20
	MCMC_indirect_write(11'd66, 68'b00001000001001001000101111000100010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd67, 68'b00001000110010010000010100000001000000101010000111100000000000000000); #20
	MCMC_indirect_write(11'd68, 68'b00000000000000000000000000000000000000000000000000000000111101011001); #20
	MCMC_indirect_write(11'd69, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd70, 68'b01101100101111011011011010011110001000011000100010110000000010011111); #20
	MCMC_indirect_write(11'd71, 68'b00010000011101110001110110001011100011100010010000001000101101000100); #20
	MCMC_indirect_write(11'd72, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd73, 68'b01011110110011001001101011101001100001111110101100000000000000000000); #20
	MCMC_indirect_write(11'd74, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd75, 68'b00011011100110001010000110000000010011111010101001100110001011001100); #20
	MCMC_indirect_write(11'd76, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd77, 68'b00011010100011010000110110101010100000000000000000000000101101100110); #20
	MCMC_indirect_write(11'd78, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd79, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd80, 68'b01100000010111101011110101000111100111011011110010110011111011011111); #20
	MCMC_indirect_write(11'd81, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd82, 68'b00111110010110000010001000001010110000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd83, 68'b00100000110011110001011001000111000001101111001011000010110000001111); #20
	MCMC_indirect_write(11'd84, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd85, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd86, 68'b00000111101110100000000101110110100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd87, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd88, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd89, 68'b00110011000001011001001100100010010010110100010000101001011101100111); #20
	MCMC_indirect_write(11'd90, 68'b00000000000000000000000000000000000000000000000000000010010011110010); #20
	MCMC_indirect_write(11'd91, 68'b00110110010110111001011010000111000100101111000011101010000111011111); #20
	MCMC_indirect_write(11'd92, 68'b01011000111011111100000100000100001010110000000011010011010001111101); #20
	MCMC_indirect_write(11'd93, 68'b01110000011101011010111111011010110110100101111100101011010000001010); #20
	MCMC_indirect_write(11'd94, 68'b01011011111010010100100110110000111000010100010010001100001100001000); #20
	MCMC_indirect_write(11'd95, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd96, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd97, 68'b10000000010110011011101101010000011001100000010111110010111010010011); #20
	MCMC_indirect_write(11'd98, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd99, 68'b01011101111010000100110000000110000111111100000101110011010000100000); #20
	MCMC_indirect_write(11'd100, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd101, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd102, 68'b10100011100011101101101111100011001001010101111100010000001100011110); #20
	MCMC_indirect_write(11'd103, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd104, 68'b00010100111110011001101111110101010100010010110100101000000101011000); #20
	MCMC_indirect_write(11'd105, 68'b00111010110100011001110110010110010010011000000111000000000000000000); #20
	MCMC_indirect_write(11'd106, 68'b00010100100111101001100000111011100001110010010010100010000111111110); #20
	MCMC_indirect_write(11'd107, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd108, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd109, 68'b00111010111001001011001100010000110100110111000010001011100101110001); #20
	MCMC_indirect_write(11'd110, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd111, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd112, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd113, 68'b00000111101101000000000000000000000000101100111100000000110010110101); #20
	MCMC_indirect_write(11'd114, 68'b00101000001001101001010100011110010010101111000101100101100110101011); #20
	MCMC_indirect_write(11'd115, 68'b00000000000000000000000000000000000001100000110000000011011111100100); #20
	MCMC_indirect_write(11'd116, 68'b00100110001101111001001000011011110000101010010000000011100011111101); #20
	MCMC_indirect_write(11'd117, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd118, 68'b00110000000110110001001011010001000001100001101010100001000010101000); #20
	MCMC_indirect_write(11'd119, 68'b00101101000001100000001010001000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd120, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd121, 68'b00000011000011101000000000000000000000010001011100000010000000001110); #20
	MCMC_indirect_write(11'd122, 68'b01110001001100100011001011111010010101101001111011101011000000100100); #20
	MCMC_indirect_write(11'd123, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd124, 68'b00101111000110001010100011010100110100010000110011101001111010001000); #20
	MCMC_indirect_write(11'd125, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd126, 68'b01010010000110010001111011100110100100010011010011001101010011111111); #20
	MCMC_indirect_write(11'd127, 68'b10111110111011011110101000111111101110110110000000110000000000000000); #20
	MCMC_indirect_write(11'd128, 68'b00010000000000000000100000000000000001000000000000000010000000000000); #20
	MCMC_indirect_write(11'd129, 68'b00001101000110111000101011000110110001000111111110000000111100001011); #20
	MCMC_indirect_write(11'd130, 68'b00100010111011001001100001001100010010111000101110000010111100101111); #20
	MCMC_indirect_write(11'd131, 68'b00010100010010010000000010101101000010011111100011100000000000000000); #20
	MCMC_indirect_write(11'd132, 68'b00110001001000110000011101111000010010001110110100000011000000101000); #20
	MCMC_indirect_write(11'd133, 68'b00011001011000110001000101011011100001100000110001100100100010000100); #20
	MCMC_indirect_write(11'd134, 68'b00000000000000000000000000000000000001100000000110100111011100000000); #20
	MCMC_indirect_write(11'd135, 68'b00010110000111101000100110110111000000011111100011100010000010101001); #20
	MCMC_indirect_write(11'd136, 68'b00101100000000000000101011000011100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd137, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd138, 68'b00000000000000000000010101101110000011000111001111100011011010101111); #20
	MCMC_indirect_write(11'd139, 68'b01100110010001111011101000110100010111011010100110101110110000010101); #20
	MCMC_indirect_write(11'd140, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd141, 68'b00110011010100100010000011000011110101001101101101001000111110101000); #20
	MCMC_indirect_write(11'd142, 68'b00000000000000000000000000000000000000101101010000000100111100010101); #20
	MCMC_indirect_write(11'd143, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd144, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd145, 68'b00010000011010100000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd146, 68'b00000000000000000000000000000000000000000000000000000001010001101001); #20
	MCMC_indirect_write(11'd147, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd148, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd149, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd150, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd151, 68'b01010001101011111001101101010111010001110010010001100000000000000000); #20
	MCMC_indirect_write(11'd152, 68'b00111101101111001010100111110000000011110001110011100111101001011110); #20
	MCMC_indirect_write(11'd153, 68'b00000000000000000000000000000000000000000000000000000011011101101000); #20
	MCMC_indirect_write(11'd154, 68'b11011010011010110110000011100110111110110101001000011100001000010111); #20
	MCMC_indirect_write(11'd155, 68'b00001001111100011000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd156, 68'b00111011001100001000101110100010100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd157, 68'b00101011111110101001011110100110000100101000001101001110000111101001); #20
	MCMC_indirect_write(11'd158, 68'b01000010011111100010101101101000110111000111000110101101000101110000); #20
	MCMC_indirect_write(11'd159, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd160, 68'b00000110110001000000110001111100100000110100000010000000000101111101); #20
	MCMC_indirect_write(11'd161, 68'b00010101001111110000000000100101010000000000000000000010010010110100); #20
	MCMC_indirect_write(11'd162, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd163, 68'b01111110001100100010110100010000110011111000001111101000011111101100); #20
	MCMC_indirect_write(11'd164, 68'b01011001011111111010000111011000100101110010110111101110000011111100); #20
	MCMC_indirect_write(11'd165, 68'b00010101111000010000100110110000100001111010010110100000001110111100); #20
	MCMC_indirect_write(11'd166, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd167, 68'b00100001001111010001011010100101010011011011100101100010111011111010); #20
	MCMC_indirect_write(11'd168, 68'b00101111110101101010010010111010010010010101110110000010010101100111); #20
	MCMC_indirect_write(11'd169, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd170, 68'b01000011001001010011100000001011000110001010011100001111100110010110); #20
	MCMC_indirect_write(11'd171, 68'b00011110101011011000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd172, 68'b01000100011001100010110011100101110101000110100010100111100000000111); #20
	MCMC_indirect_write(11'd173, 68'b00000000000000000000000110010100110001001110010111100011110011111111); #20
	MCMC_indirect_write(11'd174, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd175, 68'b00100000110000010000111100110000000000000000000000000110010000101110); #20
	MCMC_indirect_write(11'd176, 68'b01000000010001101001000011000001100010011101011101100111100001110110); #20
	MCMC_indirect_write(11'd177, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd178, 68'b00100001010010110001111010100110110100100100111001101010111011110111); #20
	MCMC_indirect_write(11'd179, 68'b00111101001101000010011010110010010101100010101110101010001010101101); #20
	MCMC_indirect_write(11'd180, 68'b00101100111011110001010001000110010000001001100010100000000000000000); #20
	MCMC_indirect_write(11'd181, 68'b00000000000000000000110101110101000001001110101010100101101100110001); #20
	MCMC_indirect_write(11'd182, 68'b10000010111001010011101111000001110111000010011000010000011111100011); #20
	MCMC_indirect_write(11'd183, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd184, 68'b00010000001101110000011001101100010001100111000011101000010110010011); #20
	MCMC_indirect_write(11'd185, 68'b00000111101010011000101001111101100001010011100110000110010111101110); #20
	MCMC_indirect_write(11'd186, 68'b00111001001011100001011000000001100000101000000111100101101100110001); #20
	MCMC_indirect_write(11'd187, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd188, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd189, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd190, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd191, 68'b00011101110100110000000000000000000010100001100001100011001011011010); #20
	MCMC_indirect_write(11'd192, 68'b00011000000000000000110000000000000001100000000000000011000000000000); #20
	MCMC_indirect_write(11'd193, 68'b00010110110000101000110110011010110001100111110110100011010000011010); #20
	MCMC_indirect_write(11'd194, 68'b00010010100111010001000100001011100010010010100000000110011011110100); #20
	MCMC_indirect_write(11'd195, 68'b00000000000000000000010110110101110010001100010100100101111100101100); #20
	MCMC_indirect_write(11'd196, 68'b00000000000000000000000000000000000000000000000000000011001010001000); #20
	MCMC_indirect_write(11'd197, 68'b00011100000011011001010001101110100001011111011100000100111110001001); #20
	MCMC_indirect_write(11'd198, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd199, 68'b01000000011110000010001010101000010010000110000101000101000110100010); #20
	MCMC_indirect_write(11'd200, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd201, 68'b00000000001001001000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd202, 68'b00110011001111010010000111010010100011111101100100101001101010100110); #20
	MCMC_indirect_write(11'd203, 68'b01000010111011000001111010110101000010000011011100100010111101000001); #20
	MCMC_indirect_write(11'd204, 68'b00100001100110110001101110100100100100110111100111100111100010111011); #20
	MCMC_indirect_write(11'd205, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd206, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd207, 68'b00010011110000010000000000000000000000111010000010000001010000001101); #20
	MCMC_indirect_write(11'd208, 68'b00101001000001001000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd209, 68'b00000011101010111000000010011111010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd210, 68'b00000000000000000000000000000000000001110000101010000101010101011100); #20
	MCMC_indirect_write(11'd211, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd212, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd213, 68'b00000000000000000000000000000000000010100111011100100000000000000000); #20
	MCMC_indirect_write(11'd214, 68'b00000010110001100000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd215, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd216, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd217, 68'b01010111010110011010011100001001100100011011011101000100101001100011); #20
	MCMC_indirect_write(11'd218, 68'b01010010001010110010111101100110110111010101111111110010011100110000); #20
	MCMC_indirect_write(11'd219, 68'b10101011100111010101100101000111001010110100100010110100000001101011); #20
	MCMC_indirect_write(11'd220, 68'b00000000000000000000011111000110100000100101011110100000001100010000); #20
	MCMC_indirect_write(11'd221, 68'b00000000000000000000010100110010100000011101000100100000000000000000); #20
	MCMC_indirect_write(11'd222, 68'b00000001001001110000010110010100110000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd223, 68'b01001111111000000010101100000001000110001001011111101110000110010110); #20
	MCMC_indirect_write(11'd224, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd225, 68'b01000100010000001001100010101101110110101110001000010010010100100000); #20
	MCMC_indirect_write(11'd226, 68'b00110000001001101011000010001001100110000111011100001110110011000001); #20
	MCMC_indirect_write(11'd227, 68'b00101110111101111010001010111011010010010011101111000011110101011010); #20
	MCMC_indirect_write(11'd228, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd229, 68'b01001001111110101000111011111111110000100000110100000100000111111110); #20
	MCMC_indirect_write(11'd230, 68'b00001110010000101001001011010010100011101101100110100110100011101111); #20
	MCMC_indirect_write(11'd231, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd232, 68'b10100001000010111110011000010111001110000100000000011011100110110111); #20
	MCMC_indirect_write(11'd233, 68'b01110110011011001011011110010111010110101111000101001111010111010011); #20
	MCMC_indirect_write(11'd234, 68'b01000111101001101010110111110000100110111010100010001011000011001100); #20
	MCMC_indirect_write(11'd235, 68'b00100011111001101000000110111000100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd236, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd237, 68'b10000111000000011011100000011110010101001111100100101100110011000010); #20
	MCMC_indirect_write(11'd238, 68'b01010001101101100010110101110011000101000101010001101111011101011101); #20
	MCMC_indirect_write(11'd239, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd240, 68'b00000000000000000000000111011011110000000000000000000000111010100001); #20
	MCMC_indirect_write(11'd241, 68'b00000000000000000000000000000000000000110010010111000001100000001100); #20
	MCMC_indirect_write(11'd242, 68'b01101111010110011011100011111100100101110111001000000110000111101110); #20
	MCMC_indirect_write(11'd243, 68'b01000001100010011000111001011011110000000000000000000010000100000011); #20
	MCMC_indirect_write(11'd244, 68'b10101100101000000100011000101011011001001100101111010000111000010110); #20
	MCMC_indirect_write(11'd245, 68'b00011010000010101001000011001111010011111010001010000011011000101000); #20
	MCMC_indirect_write(11'd246, 68'b00000001100100011000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd247, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd248, 68'b11100000010101100110111111111110001111001101101001011100000111111000); #20
	MCMC_indirect_write(11'd249, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd250, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd251, 68'b00000000000000000000011110000010000001101001111100100110000000101110); #20
	MCMC_indirect_write(11'd252, 68'b00010011001011110000100110000001010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd253, 68'b01011001010011000011110001001110000110010110000010001111101011111100); #20
	MCMC_indirect_write(11'd254, 68'b00011111011100000000000000000000000000000010111000100000000000000000); #20
	MCMC_indirect_write(11'd255, 68'b00000000000000000000000000000000000000001101101101000000000000000000); #20
	MCMC_indirect_write(11'd256, 68'b00100000000000000001000000000000000010000000000000000100000000000000); #20
	MCMC_indirect_write(11'd257, 68'b00101000100010010000111000010010010001111001001101000100011110111101); #20
	MCMC_indirect_write(11'd258, 68'b00111000000100011000111011111101000011001001111010000100011110111000); #20
	MCMC_indirect_write(11'd259, 68'b00001001111010010000011101010111000001001000001011000001000001111110); #20
	MCMC_indirect_write(11'd260, 68'b00100111111010110000011100101011100010111111011100100101110001011011); #20
	MCMC_indirect_write(11'd261, 68'b00000110010000011000000000000000000000001111010111100010100001011000); #20
	MCMC_indirect_write(11'd262, 68'b00010010001000101000111001010101110010001010100011000010110110101110); #20
	MCMC_indirect_write(11'd263, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd264, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd265, 68'b01001011000001000001101111101000010100111100100111101101100110000011); #20
	MCMC_indirect_write(11'd266, 68'b00001010010100110000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd267, 68'b00000101101011010000100100110101110000110100110001100000000000000000); #20
	MCMC_indirect_write(11'd268, 68'b01011100101101101010100111100001010100101011001100001000001001011000); #20
	MCMC_indirect_write(11'd269, 68'b01111010001110101101001111111000011001110010011011110101001100101001); #20
	MCMC_indirect_write(11'd270, 68'b01011010000000000011101100001110000111010100010000001110001100010101); #20
	MCMC_indirect_write(11'd271, 68'b01111011110100000011101101001100100111110101011101101101111001101110); #20
	MCMC_indirect_write(11'd272, 68'b01001101000010011010001110011110110100100101110011001010000110001011); #20
	MCMC_indirect_write(11'd273, 68'b01001010011101111010001011100001000011111001001100000101010100011001); #20
	MCMC_indirect_write(11'd274, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd275, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd276, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd277, 68'b00011000000000100000011010111000010001110011010010100001011011001001); #20
	MCMC_indirect_write(11'd278, 68'b01101000110100111011010010110011110101101001000010100111111110000111); #20
	MCMC_indirect_write(11'd279, 68'b00110101110100000000110100101110010010111100111110001001110100111100); #20
	MCMC_indirect_write(11'd280, 68'b00000000000000000000000000000000000001000110110101000000110100110001); #20
	MCMC_indirect_write(11'd281, 68'b00000000000000000000000000000000000000101111011101000000000000000000); #20
	MCMC_indirect_write(11'd282, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd283, 68'b00011100011011011000001001011000010000000000000000000110001011010000); #20
	MCMC_indirect_write(11'd284, 68'b00000000000000000000011110111101100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd285, 68'b00111111101000101001100110001010100101000100011110101011110111100011); #20
	MCMC_indirect_write(11'd286, 68'b00000000000000000000011010100110010010010101111100001000100001111010); #20
	MCMC_indirect_write(11'd287, 68'b01110110110101101011100111000101010111011111010011010000110111000010); #20
	MCMC_indirect_write(11'd288, 68'b11000111001111111101010111000101101000100100000010101100110100001100); #20
	MCMC_indirect_write(11'd289, 68'b00001010110101101000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd290, 68'b01110111011000001011110000001000110111110111101100010010110111000111); #20
	MCMC_indirect_write(11'd291, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd292, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd293, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd294, 68'b01001001111011100010101010111000110011000011001011100101000100011010); #20
	MCMC_indirect_write(11'd295, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd296, 68'b00000000000000000000011110110010110001110110011110100100011100110111); #20
	MCMC_indirect_write(11'd297, 68'b10010011100100111101110110000001001101010001000011111100111000000101); #20
	MCMC_indirect_write(11'd298, 68'b00011101001001110000100011001001110001101011001101000110011101100001); #20
	MCMC_indirect_write(11'd299, 68'b00110111110010111011011011111000110110101110001111101110010001100001); #20
	MCMC_indirect_write(11'd300, 68'b00000000000000000000000111000010110010000010101111000100111100011110); #20
	MCMC_indirect_write(11'd301, 68'b01000000000001000001100100001011100010100100111000100101001010001010); #20
	MCMC_indirect_write(11'd302, 68'b00111110100000111001111011100101100100101100001010001010101100111000); #20
	MCMC_indirect_write(11'd303, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd304, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd305, 68'b01011101000000010010100011011000100011001101111000000110110011010000); #20
	MCMC_indirect_write(11'd306, 68'b01010110001001101011111011101000100111111101000000101011100000110000); #20
	MCMC_indirect_write(11'd307, 68'b00011111100001100000110110111101010000010001011101000000101010001010); #20
	MCMC_indirect_write(11'd308, 68'b00101010101011111000101111101010110000101101100100100000011111100101); #20
	MCMC_indirect_write(11'd309, 68'b00101010111001011000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd310, 68'b00110001100110110010010000010000010101101010100110001110111000111011); #20
	MCMC_indirect_write(11'd311, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd312, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd313, 68'b00000000000000000000000000000000000000000000000000000000101110000101); #20
	MCMC_indirect_write(11'd314, 68'b00110100001100110001101010101101010011000001000110101000000101100110); #20
	MCMC_indirect_write(11'd315, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd316, 68'b00101010100001110001101111111100000011110001000000001010011110100110); #20
	MCMC_indirect_write(11'd317, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd318, 68'b01111010001001001010000001100011010001101101001100100001000100110010); #20
	MCMC_indirect_write(11'd319, 68'b01101111011110001011100100101000110110110100101001101110000000110001); #20
	MCMC_indirect_write(11'd320, 68'b00101000000000000001010000000000000010100000000000000101000000000000); #20
	MCMC_indirect_write(11'd321, 68'b00100001010111011001011000010000000010100111111110000101000111111000); #20
	MCMC_indirect_write(11'd322, 68'b00010000010100110000100101111111100001101101001100000000110001010100); #20
	MCMC_indirect_write(11'd323, 68'b00110100110010111001010100100011010011000100110111100010011011001010); #20
	MCMC_indirect_write(11'd324, 68'b00000000000000000000000000000000000010110001100101000110001101011011); #20
	MCMC_indirect_write(11'd325, 68'b00010000000010000001010110100011010110010100110011101110011110011101); #20
	MCMC_indirect_write(11'd326, 68'b00011001011000000001101010110100110011010111110011100110000100100010); #20
	MCMC_indirect_write(11'd327, 68'b00000000000000000000111111010010000100000011001110000111000100101111); #20
	MCMC_indirect_write(11'd328, 68'b10100111101001100100001010100000101000110110000101001011011100001111); #20
	MCMC_indirect_write(11'd329, 68'b01010101100010010011000101100100110101101101011001101101000101010001); #20
	MCMC_indirect_write(11'd330, 68'b01010001111100000010001101001011010101100100101111001101110010100111); #20
	MCMC_indirect_write(11'd331, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd332, 68'b01101010110100001010110010000110000101100110011111101100010110110010); #20
	MCMC_indirect_write(11'd333, 68'b00001100001110000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd334, 68'b00100111010110111000011101110100000000000000000000000011111101011011); #20
	MCMC_indirect_write(11'd335, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd336, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd337, 68'b10011111100101000110011000000010011010110110111100010101011101100000); #20
	MCMC_indirect_write(11'd338, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd339, 68'b00111011110101010010010101010101110100011010100010101100101001100101); #20
	MCMC_indirect_write(11'd340, 68'b00001111111100000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd341, 68'b01000010011010010000110100110111010011000110000010000001011101010111); #20
	MCMC_indirect_write(11'd342, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd343, 68'b01000000100010101010000101011100100100101010001001101001011101101001); #20
	MCMC_indirect_write(11'd344, 68'b01000110010000101001101011010011000000111000000011100000000000000000); #20
	MCMC_indirect_write(11'd345, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd346, 68'b01110100111010110010101111110011010110000001110000101011011110011000); #20
	MCMC_indirect_write(11'd347, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd348, 68'b01010000111001000011011000010110110110011001000011101101000100110011); #20
	MCMC_indirect_write(11'd349, 68'b00000000000000000000000000000000000000000000000000000100000000100011); #20
	MCMC_indirect_write(11'd350, 68'b00010101101010011001010111010001000001111000001110000000000000000000); #20
	MCMC_indirect_write(11'd351, 68'b10001100111010111100011001011111001001000100001011001101001101011001); #20
	MCMC_indirect_write(11'd352, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd353, 68'b00100111010001001000000000101010100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd354, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd355, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd356, 68'b00100100010101111000001010010001110001000011001110000101010000100111); #20
	MCMC_indirect_write(11'd357, 68'b00010001100101111000111111011001010010110000111110100010111011111010); #20
	MCMC_indirect_write(11'd358, 68'b00100001000111100000000000000000000000101011111100000000000000000000); #20
	MCMC_indirect_write(11'd359, 68'b01000001101000101010010011000010110100011010110100000110100110000001); #20
	MCMC_indirect_write(11'd360, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd361, 68'b10100100010101001100101010101000101000001111000001010000100101001110); #20
	MCMC_indirect_write(11'd362, 68'b10101000101000101101111011110100001011001111110011110100110010100111); #20
	MCMC_indirect_write(11'd363, 68'b10111000111110101101011110101010001100001110100111010100001010111011); #20
	MCMC_indirect_write(11'd364, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd365, 68'b10011100111011010101010101011001111010110000001000010010010000010100); #20
	MCMC_indirect_write(11'd366, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd367, 68'b01111101010100110011001110110010010101010100101000101000000101111111); #20
	MCMC_indirect_write(11'd368, 68'b01110100100001010010100110011000110110111110000101001111000001111111); #20
	MCMC_indirect_write(11'd369, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd370, 68'b00001000100111110000100001000010000000000101111010100000000000000000); #20
	MCMC_indirect_write(11'd371, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd372, 68'b01111001010100010011011010101100010111100001101011001110011011100011); #20
	MCMC_indirect_write(11'd373, 68'b00000000000000000000000000000000000000000000000000000100000000000010); #20
	MCMC_indirect_write(11'd374, 68'b10011101110111110100001110010011010110110110011010001110001110010101); #20
	MCMC_indirect_write(11'd375, 68'b00000101000111010000010010101111010001100010000101000000000000000000); #20
	MCMC_indirect_write(11'd376, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd377, 68'b10110101101010011110001000000010111011000110000000110001000110100111); #20
	MCMC_indirect_write(11'd378, 68'b01011010011000000010111111011101010011101100110011000101100011001001); #20
	MCMC_indirect_write(11'd379, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd380, 68'b00010111101110010000000000000000000000000000000000000010101100111001); #20
	MCMC_indirect_write(11'd381, 68'b01011100000101010010001110100011110010000000011100001000010100010011); #20
	MCMC_indirect_write(11'd382, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd383, 68'b00011110101001000001001000010010010100010011101110001000011001010011); #20
	MCMC_indirect_write(11'd384, 68'b00110000000000000001100000000000000011000000000000000110000000000000); #20
	MCMC_indirect_write(11'd385, 68'b00101000010001001001011000110110010011010010101100000101010110000111); #20
	MCMC_indirect_write(11'd386, 68'b01001100110010100001101100110110110010001001001000000101101001101101); #20
	MCMC_indirect_write(11'd387, 68'b00001001010100011001010101010100010000111000111011100001101000110110); #20
	MCMC_indirect_write(11'd388, 68'b00101100100000010001110111111100000100101010100010001010110000011110); #20
	MCMC_indirect_write(11'd389, 68'b01100101011010000010100100010010000100100011100011100101111110011101); #20
	MCMC_indirect_write(11'd390, 68'b00110111111101101000010111101011110000100011010001100000000000000000); #20
	MCMC_indirect_write(11'd391, 68'b01000101011100001001111101110100100010111110001001000001000101100001); #20
	MCMC_indirect_write(11'd392, 68'b00110011000111110010001011010000010011010100010000000101101110001010); #20
	MCMC_indirect_write(11'd393, 68'b01110000111000011011011110101111110011101101000011101100101001101000); #20
	MCMC_indirect_write(11'd394, 68'b00111111100010000010001010100000000011101010011001101001011000000100); #20
	MCMC_indirect_write(11'd395, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd396, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd397, 68'b01000101100101110010100101101000110110100100000011101110111010111111); #20
	MCMC_indirect_write(11'd398, 68'b01110000010100001101011100100111011000110100110110010001100000111111); #20
	MCMC_indirect_write(11'd399, 68'b00000100010100011000101011110101110000000000000000000000110011101111); #20
	MCMC_indirect_write(11'd400, 68'b01000100110000000010010111100011110100100101101000100101011011100010); #20
	MCMC_indirect_write(11'd401, 68'b00000011100011001000101010000010100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd402, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd403, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd404, 68'b00000110001011111000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd405, 68'b00010111100001001001000010011010000011001000011110100001011100010000); #20
	MCMC_indirect_write(11'd406, 68'b00100110001010101001100100100010110101001011101111001000101011010001); #20
	MCMC_indirect_write(11'd407, 68'b00110111111111010001111100000010000100111001011011101100101111101101); #20
	MCMC_indirect_write(11'd408, 68'b10001011001100010011111101100111100111101110000110101110111101000010); #20
	MCMC_indirect_write(11'd409, 68'b10100001111010010011111011110110110111101010101001110010001111101101); #20
	MCMC_indirect_write(11'd410, 68'b00111110011111001001101011011010010111000100100110101100101110010001); #20
	MCMC_indirect_write(11'd411, 68'b01000101001001010001001010000000100010100101101101101001001100101100); #20
	MCMC_indirect_write(11'd412, 68'b00111100001000000010100110100010000111011001000110001101111001101010); #20
	MCMC_indirect_write(11'd413, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd414, 68'b00000000000000000000000000000000000000000000000000000001100101000011); #20
	MCMC_indirect_write(11'd415, 68'b10010101101110001100001011011001000111001111010100010011000001001110); #20
	MCMC_indirect_write(11'd416, 68'b01011000010101001011100111001010000101011000101100101000011011001001); #20
	MCMC_indirect_write(11'd417, 68'b10001000000001011100001000010101010110101010001001101111011010010001); #20
	MCMC_indirect_write(11'd418, 68'b00000000000000000000000000101110000001000100111100100100011101100101); #20
	MCMC_indirect_write(11'd419, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd420, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd421, 68'b01000111111001011010000000101010100100000100110100100111010111110010); #20
	MCMC_indirect_write(11'd422, 68'b01100111100001011011000010100001011000010110110110110000010001110001); #20
	MCMC_indirect_write(11'd423, 68'b00000000000000000000000000000000000000000000000000000010000010101101); #20
	MCMC_indirect_write(11'd424, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd425, 68'b01000010100110101011000101111101100100111110111010101100010110001001); #20
	MCMC_indirect_write(11'd426, 68'b00000000000000000001011101111101010000000000000000000001111011010101); #20
	MCMC_indirect_write(11'd427, 68'b01001000001001110001001111000100000011110111101100100111001110101110); #20
	MCMC_indirect_write(11'd428, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd429, 68'b01000001011111101010001110100011010010100110001001000001101010011001); #20
	MCMC_indirect_write(11'd430, 68'b00000011100100100000010011011010100010010000000101100101000001011001); #20
	MCMC_indirect_write(11'd431, 68'b00011001111110001000100101010111100010100011000110001001001101111101); #20
	MCMC_indirect_write(11'd432, 68'b01101011011010000011111100100111100111010011010001101101100000010001); #20
	MCMC_indirect_write(11'd433, 68'b00101110111111101010011000110110010101111001111011101110001011010010); #20
	MCMC_indirect_write(11'd434, 68'b10001101010011001110011000000010111100001001111111111000100000010011); #20
	MCMC_indirect_write(11'd435, 68'b00101101101101100001010010010110010010001001110101100111111001000110); #20
	MCMC_indirect_write(11'd436, 68'b01011111101110001010101101111010100110011100110110101100100111111001); #20
	MCMC_indirect_write(11'd437, 68'b01011011000010110011001101000110100110101101110111010000110101101000); #20
	MCMC_indirect_write(11'd438, 68'b01111101000011111011100011001110001000110101011100101111100111011011); #20
	MCMC_indirect_write(11'd439, 68'b01110011111010001010111100101110000110011010111111101101111111000000); #20
	MCMC_indirect_write(11'd440, 68'b01100011001010110010110111010010000110111101010011101010101010010011); #20
	MCMC_indirect_write(11'd441, 68'b00110000111110101010010001100010110101000010001110101000100010110110); #20
	MCMC_indirect_write(11'd442, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd443, 68'b01011101101010111010000001010110100101110110001000100111010011010010); #20
	MCMC_indirect_write(11'd444, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd445, 68'b01000100100110001001000000011100010001011110100011100101001000001011); #20
	MCMC_indirect_write(11'd446, 68'b00001000101011110000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd447, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd448, 68'b00111000000000000001110000000000000011100000000000000111000000000000); #20
	MCMC_indirect_write(11'd449, 68'b01000000000111001010000100011011010011100110011001100111101101101000); #20
	MCMC_indirect_write(11'd450, 68'b01000111010011010010011001011001100011000001011010000110101110010101); #20
	MCMC_indirect_write(11'd451, 68'b00101000111111110001110110110001000011010000110111000101011000000111); #20
	MCMC_indirect_write(11'd452, 68'b00110001101100111001110111101000100011101001001100000111001100000100); #20
	MCMC_indirect_write(11'd453, 68'b00011011110000010001011100101010010010100001001100000110001000100011); #20
	MCMC_indirect_write(11'd454, 68'b00010111000011101000000000000000000001010011101001000000111110110000); #20
	MCMC_indirect_write(11'd455, 68'b10000111001011101100101010100110100110111111110010100111100011011101); #20
	MCMC_indirect_write(11'd456, 68'b10000000000100101100100011101110101100100000101111110100010000010111); #20
	MCMC_indirect_write(11'd457, 68'b00111110101111010001110111000110010110000011010100101000110000001110); #20
	MCMC_indirect_write(11'd458, 68'b00110010100011000010010010010110100101100000100111101000011111101110); #20
	MCMC_indirect_write(11'd459, 68'b01001110001000000010100101100111000100001110110000101011001011010011); #20
	MCMC_indirect_write(11'd460, 68'b00110111001000110001111110010100110010001010011011000100010000110010); #20
	MCMC_indirect_write(11'd461, 68'b01001111011111011010101010110001010101110111000110000100011111001010); #20
	MCMC_indirect_write(11'd462, 68'b01101000111000001100000110101000100110100010000101001000100100111000); #20
	MCMC_indirect_write(11'd463, 68'b00101100000001101000111011100011100011111110101110000101011000011111); #20
	MCMC_indirect_write(11'd464, 68'b10101110010101000100001110001101000111101010111001101110000010011000); #20
	MCMC_indirect_write(11'd465, 68'b01010000101110000000111101111011110001000101001000000101010111000011); #20
	MCMC_indirect_write(11'd466, 68'b10001001011101000101001101011001111101001101010100010100001000011100); #20
	MCMC_indirect_write(11'd467, 68'b10101000110011111110000010100000011101100101000100111010001110110110); #20
	MCMC_indirect_write(11'd468, 68'b01010100011001100001011110001011010010101000011110100000101001010000); #20
	MCMC_indirect_write(11'd469, 68'b01100100000000101011010111001011001000011011000101001110011011011010); #20
	MCMC_indirect_write(11'd470, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd471, 68'b01001011100001100010011100010111000011011001011101100101011001101111); #20
	MCMC_indirect_write(11'd472, 68'b01000101110011010010100010011001110100110101001111100111011010001000); #20
	MCMC_indirect_write(11'd473, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd474, 68'b01101111101101010101000000001010001001010101100011110110100100011111); #20
	MCMC_indirect_write(11'd475, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd476, 68'b01101000100100101011110101011010001000111101001011110010101001010011); #20
	MCMC_indirect_write(11'd477, 68'b10001100011100001101011010110110111001000110001010110010000101010011); #20
	MCMC_indirect_write(11'd478, 68'b01001111101001101010110011010100100101011010011110001011111111111000); #20
	MCMC_indirect_write(11'd479, 68'b01001011101001111011100000110011010111100001010001001100001100000100); #20
	MCMC_indirect_write(11'd480, 68'b00000000000000000000000100100110000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd481, 68'b00110000111111101001011110011111100001011011100010000010111011001101); #20
	MCMC_indirect_write(11'd482, 68'b00000000000000000000000000000000000000000000000000000000110111111101); #20
	MCMC_indirect_write(11'd483, 68'b01100100011001100011001010101110110110001101011010001010111101111000); #20
	MCMC_indirect_write(11'd484, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd485, 68'b00110111010001100010111100000100000110100100101001101011111011100010); #20
	MCMC_indirect_write(11'd486, 68'b00111100111100010010011010010000000010011010100000100101110111110111); #20
	MCMC_indirect_write(11'd487, 68'b00010011011100011000000001101110110000000000000000000011001000110110); #20
	MCMC_indirect_write(11'd488, 68'b01100010001100010001010110010000010000001100011111000001001101111011); #20
	MCMC_indirect_write(11'd489, 68'b00010110001000101000010010110001110001110000011100000100110100001010); #20
	MCMC_indirect_write(11'd490, 68'b01011101110110111010110101000110110111001010001011000111011011000010); #20
	MCMC_indirect_write(11'd491, 68'b01001101101111010011101011101101010111011100001100101111001000101010); #20
	MCMC_indirect_write(11'd492, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd493, 68'b01011101101010011011100110101111100101110100010101001100011010110110); #20
	MCMC_indirect_write(11'd494, 68'b01101011111100110010001000001001100110000010010010001110001000101000); #20
	MCMC_indirect_write(11'd495, 68'b00101001101010100000101110101100110010101000111100000101100111000110); #20
	MCMC_indirect_write(11'd496, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd497, 68'b10010000011011011100110010111111010110001101100111001011000100001011); #20
	MCMC_indirect_write(11'd498, 68'b00011110010101001000110000000011110000000000000000000010001001100101); #20
	MCMC_indirect_write(11'd499, 68'b01001111111010000001101010000101010100111101100010100101111111100111); #20
	MCMC_indirect_write(11'd500, 68'b00111010000000000001100100100110000001001111010011000011001000101101); #20
	MCMC_indirect_write(11'd501, 68'b01001101011000101001010100100000010100011010100110000110001011110001); #20
	MCMC_indirect_write(11'd502, 68'b00010100011001001000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd503, 68'b10001111101100110011111011110010110110000101010010001000111010011011); #20
	MCMC_indirect_write(11'd504, 68'b01101110001100111011101101110110000100111111010011100110100110110110); #20
	MCMC_indirect_write(11'd505, 68'b01000101000011011010010011110010110011001110100101100111000001010111); #20
	MCMC_indirect_write(11'd506, 68'b10001100010010101100011101010110100110000111100011010010101001101100); #20
	MCMC_indirect_write(11'd507, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd508, 68'b01110110001000100100001100011110111001100010000101110100010110110101); #20
	MCMC_indirect_write(11'd509, 68'b01001100100000011010011000011010100011111110101101100101101011100111); #20
	MCMC_indirect_write(11'd510, 68'b00101111000111111001000001001001010011000000101000001000111100000010); #20
	MCMC_indirect_write(11'd511, 68'b00111111010010101000111001010100010000011110010101100000100001101101); #20
	MCMC_indirect_write(11'd512, 68'b01000000000000000010000000000000000100000000000000001000000000000000); #20
	MCMC_indirect_write(11'd513, 68'b00111011000010001010000011111000100100001110100111000111001011110011); #20
	MCMC_indirect_write(11'd514, 68'b00101110010111111001101011100100010100101001111100001001100010011101); #20
	MCMC_indirect_write(11'd515, 68'b00110010100101001010001100011000010100100000101001000100110100000100); #20
	MCMC_indirect_write(11'd516, 68'b01100001100100100010110010101110000011101001001101001000110111110100); #20
	MCMC_indirect_write(11'd517, 68'b00110001100011000000111001101000010000001011001100100001110101001000); #20
	MCMC_indirect_write(11'd518, 68'b00111001011110110001011101110011100011011010100011100110100101001001); #20
	MCMC_indirect_write(11'd519, 68'b10001010000001110101110011100111101001101011000100010000111000100101); #20
	MCMC_indirect_write(11'd520, 68'b00000000000000000000000000000000000000000000000000000001001000100010); #20
	MCMC_indirect_write(11'd521, 68'b00100100101100100001100110110000000100011101100011000011010011110001); #20
	MCMC_indirect_write(11'd522, 68'b01010110110111000001101101001100100100001100001001001101010101010100); #20
	MCMC_indirect_write(11'd523, 68'b00011011101010010001011111001000010011001111100010101001110111101000); #20
	MCMC_indirect_write(11'd524, 68'b10100010001100011100111000110001111100000011001001010011101001100000); #20
	MCMC_indirect_write(11'd525, 68'b00111101100110110010001110100100010110000010110010100101101001001010); #20
	MCMC_indirect_write(11'd526, 68'b01000001110001100010110000011011000101011100010001101100011100111001); #20
	MCMC_indirect_write(11'd527, 68'b01101010011101110010101100001101011000111011001110101111011011001111); #20
	MCMC_indirect_write(11'd528, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd529, 68'b10101000100010111100110110110000111011111111011100011000001010000110); #20
	MCMC_indirect_write(11'd530, 68'b00011011111110110000110010001011110001100100000100100100110010100100); #20
	MCMC_indirect_write(11'd531, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd532, 68'b10010011010000000100001100101010100110110001100011001001100001111110); #20
	MCMC_indirect_write(11'd533, 68'b00111000111000011001110111100111000011101000011001101001100111110101); #20
	MCMC_indirect_write(11'd534, 68'b01011111000101011011000000111111110110110001101000001100100100100101); #20
	MCMC_indirect_write(11'd535, 68'b01101101111010010100100001010100000110000001000010110011101101101100); #20
	MCMC_indirect_write(11'd536, 68'b00000000000000000001010100001001010011010001101100100111011110000101); #20
	MCMC_indirect_write(11'd537, 68'b10011001101111101101001110010011111011010000111000011000000100101000); #20
	MCMC_indirect_write(11'd538, 68'b00101001010110011000111001001000000000000000000000000000101111101110); #20
	MCMC_indirect_write(11'd539, 68'b10101010100110100101100011101010101100011010110000110100100001110100); #20
	MCMC_indirect_write(11'd540, 68'b00110001011011101000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd541, 68'b00101011011110101000011100101011100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd542, 68'b00101101110000011001100010100110000011100111011110101001100100101101); #20
	MCMC_indirect_write(11'd543, 68'b01010101011101111010001001010111100011101010110101101000010111000101); #20
	MCMC_indirect_write(11'd544, 68'b00000000000000000000000100100000010000011010110011000001011111010110); #20
	MCMC_indirect_write(11'd545, 68'b00010100111001111000010000100001000001101001011010001000100001011110); #20
	MCMC_indirect_write(11'd546, 68'b00000000000000000000001100001111000000101011000111000011111110101111); #20
	MCMC_indirect_write(11'd547, 68'b01101111001101100011101111011011000111011101110111010011010100111101); #20
	MCMC_indirect_write(11'd548, 68'b01010000000111101011111011010010100111011011101010010000110000001011); #20
	MCMC_indirect_write(11'd549, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd550, 68'b00100100110010100001100010101100000010001011101011000011111000111000); #20
	MCMC_indirect_write(11'd551, 68'b00101000100001110001011000001111010011000110111100101011010001011110); #20
	MCMC_indirect_write(11'd552, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd553, 68'b00101100100101100000000111111001010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd554, 68'b10011000111000101101001011001001011010110101001100110111111001101110); #20
	MCMC_indirect_write(11'd555, 68'b00000000100111001000110101110011000010001100101001000100111101000101); #20
	MCMC_indirect_write(11'd556, 68'b10001000110110101101011010111101111011001110100100111100011100101001); #20
	MCMC_indirect_write(11'd557, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd558, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd559, 68'b01011010100100111010111000100110010100101000111101101100110100110100); #20
	MCMC_indirect_write(11'd560, 68'b01010100011010100001111010010110010010100010011111100010011011011111); #20
	MCMC_indirect_write(11'd561, 68'b10000011000111111011110000000010001000001000101101001100101000101111); #20
	MCMC_indirect_write(11'd562, 68'b10100010101101011100111100011101001000011001100110010000011000110111); #20
	MCMC_indirect_write(11'd563, 68'b01010101101111010010110111001111110101001111000010101001010010111001); #20
	MCMC_indirect_write(11'd564, 68'b10000100111010001011100110011000000111001010100110001100110101010010); #20
	MCMC_indirect_write(11'd565, 68'b00101110000000011010001111110001110011000100101111100100011001000101); #20
	MCMC_indirect_write(11'd566, 68'b01101111100100010011111110010110000110001111100111001110000011111101); #20
	MCMC_indirect_write(11'd567, 68'b00000000000000000000000000000000000000000000000000000010110111010011); #20
	MCMC_indirect_write(11'd568, 68'b01001111001001011010111100011110110110000111111001110000011111111010); #20
	MCMC_indirect_write(11'd569, 68'b10011000100101011011110111010000011001110010001110010010011110010000); #20
	MCMC_indirect_write(11'd570, 68'b00111111000111011010000100101000110100001101110011100100100111110101); #20
	MCMC_indirect_write(11'd571, 68'b00110010001000001001000110000110000011111111101000100111001101111011); #20
	MCMC_indirect_write(11'd572, 68'b00111001100000100001010101101001000011111101101110000110011000000010); #20
	MCMC_indirect_write(11'd573, 68'b10100001100101000101011100010111101100110101101010011011010101110010); #20
	MCMC_indirect_write(11'd574, 68'b01011111111101100100010110011001111000000001011100101010110100110111); #20
	MCMC_indirect_write(11'd575, 68'b00000100010111010000101010100010110011001010010011100011000101101011); #20
	MCMC_indirect_write(11'd576, 68'b01001000000000000010010000000000000100100000000000001001000000000000); #20
	MCMC_indirect_write(11'd577, 68'b01000110100000001010010001111011110100011101010111101010010000111101); #20
	MCMC_indirect_write(11'd578, 68'b01010010010101001010000101010101010101101010010000000110101101011011); #20
	MCMC_indirect_write(11'd579, 68'b00100001010101001001001101110110110011101010010000001010110100010000); #20
	MCMC_indirect_write(11'd580, 68'b01011110011011110011001101100110110110111010011111001101111111110010); #20
	MCMC_indirect_write(11'd581, 68'b00110011000100111001101000101010010101100111001001001001110001101000); #20
	MCMC_indirect_write(11'd582, 68'b01100100101010001011010001100001010110000111100100001110000111001100); #20
	MCMC_indirect_write(11'd583, 68'b10001100011101001100110101101010101010001100111110010010110111100100); #20
	MCMC_indirect_write(11'd584, 68'b01101111111011101010100110100011000100000110101001101001000011011001); #20
	MCMC_indirect_write(11'd585, 68'b10001101111001101011111110011101100011101010010000101011111010111101); #20
	MCMC_indirect_write(11'd586, 68'b01110000110100000011000010001011110110110111110001101110100011110000); #20
	MCMC_indirect_write(11'd587, 68'b00000000000000000000000101101110100010100001001000100100101001010001); #20
	MCMC_indirect_write(11'd588, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd589, 68'b11101010101011001111011110101001101101110110010100011110111010101110); #20
	MCMC_indirect_write(11'd590, 68'b10110101010100100101100100111111011100001011111011110110101111011100); #20
	MCMC_indirect_write(11'd591, 68'b01011000110011001001110011110110110011110111010010000101111000001100); #20
	MCMC_indirect_write(11'd592, 68'b00001100001000010000000100000111000000001010011001000000000000000000); #20
	MCMC_indirect_write(11'd593, 68'b00011101010111101000010111110001000000010001000011000000000000000000); #20
	MCMC_indirect_write(11'd594, 68'b00101001010010111001010011000010000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd595, 68'b00010000110010001001001110101100000001011011101010100111000111011010); #20
	MCMC_indirect_write(11'd596, 68'b00010110000100110000101011011011100101011011010010101111010001010000); #20
	MCMC_indirect_write(11'd597, 68'b00001100010000110000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd598, 68'b00110110011101010011010101011101010101111100010001101110101001011000); #20
	MCMC_indirect_write(11'd599, 68'b00111011101011001010001110010011000011001111101000100100001000110111); #20
	MCMC_indirect_write(11'd600, 68'b01000110111111100010000111110000010110000111110010000100110001011110); #20
	MCMC_indirect_write(11'd601, 68'b01110000100110000100000101101101001010010110110000110111110010000110); #20
	MCMC_indirect_write(11'd602, 68'b01111010100011111011110000100101011001001010101111101111000110011111); #20
	MCMC_indirect_write(11'd603, 68'b01100111010010000010110111111010010010101110011010000100101010101101); #20
	MCMC_indirect_write(11'd604, 68'b01110001110011101011101111000000101000111011100111010011010001011011); #20
	MCMC_indirect_write(11'd605, 68'b00001110100001100001000000010100000011000001011111000111100101110110); #20
	MCMC_indirect_write(11'd606, 68'b00110010011110000001000010011011010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd607, 68'b11001110001100100110010100101010101100001000011101111010011110110001); #20
	MCMC_indirect_write(11'd608, 68'b11011111010111001111001010111100001010111001111010110110100011010001); #20
	MCMC_indirect_write(11'd609, 68'b00010100110010011000110111110100000000100111000111000110000110110001); #20
	MCMC_indirect_write(11'd610, 68'b00000000000000000000000000000000000000110111111001100001011010001111); #20
	MCMC_indirect_write(11'd611, 68'b01010010000100111000101010111011010001010101010110100010011011011001); #20
	MCMC_indirect_write(11'd612, 68'b00001100010000011000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd613, 68'b00000000000000000000000000000000000000000000000000000001001101100101); #20
	MCMC_indirect_write(11'd614, 68'b00011111100101010001100000010000010001100100110001100000000000000000); #20
	MCMC_indirect_write(11'd615, 68'b00110010011001011000011010010110010000010011010010100010011010010010); #20
	MCMC_indirect_write(11'd616, 68'b00000000000000000001000000001001010001000010101011000100011110111111); #20
	MCMC_indirect_write(11'd617, 68'b01011100010000000001010010110011000011011010111011100100101011011110); #20
	MCMC_indirect_write(11'd618, 68'b01100100110001010011000001111110100111001010100010001110001111101011); #20
	MCMC_indirect_write(11'd619, 68'b01000001001101111001100111001000000110101010001100101111000011101100); #20
	MCMC_indirect_write(11'd620, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd621, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd622, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd623, 68'b10000010001010000010011011011010010101010010011110000101110100100000); #20
	MCMC_indirect_write(11'd624, 68'b00111000101000110010111010111001110100000110110100001011001110001001); #20
	MCMC_indirect_write(11'd625, 68'b00010001011110000001001110011110000011101011011001000111000001101100); #20
	MCMC_indirect_write(11'd626, 68'b00111110010011111010101111000010100100101000010000001001010011001111); #20
	MCMC_indirect_write(11'd627, 68'b00111100111001101010110101001100000110010011000101001001100010000001); #20
	MCMC_indirect_write(11'd628, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd629, 68'b01010111101101110010001001011010010100000110010001101100011011111110); #20
	MCMC_indirect_write(11'd630, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd631, 68'b01011100001100001001111111111001100011110111000011100011000001000000); #20
	MCMC_indirect_write(11'd632, 68'b10011111100000101110000001000100001100111000111001011011010111101000); #20
	MCMC_indirect_write(11'd633, 68'b00000000000000000000111111101110110000100011001100000000000000000000); #20
	MCMC_indirect_write(11'd634, 68'b00011011001110001000000011000101110000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd635, 68'b00110000010110001000101000001001110000000001101110100001010001101001); #20
	MCMC_indirect_write(11'd636, 68'b11001100011010111101010111111011111001011000000000110111101010001001); #20
	MCMC_indirect_write(11'd637, 68'b01011000000111111011000111001110100110100011110110001011001101011100); #20
	MCMC_indirect_write(11'd638, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd639, 68'b01101010000111110100000011111011100111001101011001001101110011001101); #20
	MCMC_indirect_write(11'd640, 68'b01010000000000000010100000000000000101000000000000001010000000000000); #20
	MCMC_indirect_write(11'd641, 68'b01000111100000011010011001001001000101111010001000101010101001011001); #20
	MCMC_indirect_write(11'd642, 68'b01101001000101001011000111101010100100001001000101101011000100101101); #20
	MCMC_indirect_write(11'd643, 68'b01001011000100101010100010011000000101000011010100010001000111011011); #20
	MCMC_indirect_write(11'd644, 68'b01010100110011011011110010111011000101110000110000001010110110001000); #20
	MCMC_indirect_write(11'd645, 68'b01010100110111000011010011100101110100100101001000101100100010001010); #20
	MCMC_indirect_write(11'd646, 68'b01100010011011001011111101100000010111010001010010101111100011111000); #20
	MCMC_indirect_write(11'd647, 68'b00110011000100100001101101111101010001010111101101000011000101111110); #20
	MCMC_indirect_write(11'd648, 68'b01000011101111101010010011101100000100100001001001001011110101111100); #20
	MCMC_indirect_write(11'd649, 68'b00111000100110000001110010011111100011000111110010101010011101101100); #20
	MCMC_indirect_write(11'd650, 68'b00010100001100010000011110011101100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd651, 68'b11000001100110110110001010110010111011110101101101110111110011111011); #20
	MCMC_indirect_write(11'd652, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd653, 68'b10000000100011010101000011111110101000101101010111101111110111101000); #20
	MCMC_indirect_write(11'd654, 68'b01101110110000000011011001111010010111010011000101010000011001010111); #20
	MCMC_indirect_write(11'd655, 68'b10111111111101101101011101010111101011001100001101101110001110100010); #20
	MCMC_indirect_write(11'd656, 68'b01110100011111110010111010101010000110000010101001001010101100000001); #20
	MCMC_indirect_write(11'd657, 68'b10001010101001010011011111001110100110010111100100001011111100000110); #20
	MCMC_indirect_write(11'd658, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd659, 68'b00010000010110110000010010101001110010010101010111000110010010011001); #20
	MCMC_indirect_write(11'd660, 68'b01000000000100111010000001001111100010110001110011100011011110110000); #20
	MCMC_indirect_write(11'd661, 68'b10011011110001011101001000011101001000110111111101110011011101111110); #20
	MCMC_indirect_write(11'd662, 68'b10010001100011100100000110110110110111010001111011110101110000000100); #20
	MCMC_indirect_write(11'd663, 68'b01001101111101100011101011111001011000111111001000010110110000001110); #20
	MCMC_indirect_write(11'd664, 68'b00100110011101110001100010001011110101101111011001001101001111100101); #20
	MCMC_indirect_write(11'd665, 68'b10000110010001000101111110001001011111100001100011111101010101110011); #20
	MCMC_indirect_write(11'd666, 68'b00001100010111010010001110100101110100100001011010001101000100100111); #20
	MCMC_indirect_write(11'd667, 68'b10001100001001000101100000010101011010101111110111110110011111101111); #20
	MCMC_indirect_write(11'd668, 68'b01000011110111100010100100100010100100001001010011001100110110000001); #20
	MCMC_indirect_write(11'd669, 68'b10111010011101001110011011110011001011000001011101110111000111010000); #20
	MCMC_indirect_write(11'd670, 68'b01011010000100110011011011010011100110101010101100001000011001010011); #20
	MCMC_indirect_write(11'd671, 68'b00111011011011110010000011100110100100100001101110001000010001001011); #20
	MCMC_indirect_write(11'd672, 68'b00001010000101101000101010110000000011001111000010101000100101000011); #20
	MCMC_indirect_write(11'd673, 68'b00111001000011100001011000110111100011110000010010100010101011001001); #20
	MCMC_indirect_write(11'd674, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd675, 68'b01001110001100010001110000001100000100001100001010001001000011110100); #20
	MCMC_indirect_write(11'd676, 68'b10001101010100000100011100100101101010110001110110110011001000001010); #20
	MCMC_indirect_write(11'd677, 68'b01110111100101001100010000001111001000100000011111010111110000000001); #20
	MCMC_indirect_write(11'd678, 68'b00100101010001011001001001011100010010101011110001000101101100101111); #20
	MCMC_indirect_write(11'd679, 68'b01000110010111111001101101111110100011010111010011101000001000111001); #20
	MCMC_indirect_write(11'd680, 68'b01111100011011001100000011110000001100000010100100111000111111011110); #20
	MCMC_indirect_write(11'd681, 68'b10011111001101111011110111110000110101001111110011001011111110111010); #20
	MCMC_indirect_write(11'd682, 68'b00110101010110000000110001111111100001101011111011100101100001111010); #20
	MCMC_indirect_write(11'd683, 68'b01001100110010000000110000001000000001011111001011100011000100001100); #20
	MCMC_indirect_write(11'd684, 68'b01101110000110010010110010111010100101000110010111101101101011011101); #20
	MCMC_indirect_write(11'd685, 68'b10101100100111111100101010101001000111110001011100101011010110011001); #20
	MCMC_indirect_write(11'd686, 68'b00011111000001010000011111111011100000111110111011000001000100110001); #20
	MCMC_indirect_write(11'd687, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd688, 68'b10001110010100011101000000001101101011001011100101111000100111011010); #20
	MCMC_indirect_write(11'd689, 68'b01011000101001001010000101011110010100101101100010100101100001001010); #20
	MCMC_indirect_write(11'd690, 68'b11011101001101110111001000000001101111101110110001111111001111000111); #20
	MCMC_indirect_write(11'd691, 68'b11011110000101001110001110001000011101010010110010111000100100010001); #20
	MCMC_indirect_write(11'd692, 68'b00111001111010010001101100111000100000110011011111000101001011101010); #20
	MCMC_indirect_write(11'd693, 68'b00101000001101101010011000111111010100110110010100001010111100100010); #20
	MCMC_indirect_write(11'd694, 68'b01001001100010000001010001101100010110101100011000100111010001000010); #20
	MCMC_indirect_write(11'd695, 68'b01101010101000101101000100000001011010011110101111010111000000010000); #20
	MCMC_indirect_write(11'd696, 68'b10100111010010001100111010011001111010010100110111010001011001011001); #20
	MCMC_indirect_write(11'd697, 68'b00111011111110001001110001010011110100111101001101100111110010000001); #20
	MCMC_indirect_write(11'd698, 68'b00110000010110110010100100011010110011101011010000000101111101011010); #20
	MCMC_indirect_write(11'd699, 68'b10100110110110011100100001110101010111110110000011101100110011101000); #20
	MCMC_indirect_write(11'd700, 68'b10011110000110111100001010110100001010100001111101110110100100100011); #20
	MCMC_indirect_write(11'd701, 68'b00100011001100000001110101000101000101111001111111000110101000000001); #20
	MCMC_indirect_write(11'd702, 68'b01100101010001101010001110011110000011001010101000100111100010000000); #20
	MCMC_indirect_write(11'd703, 68'b10100100000111101110101100111111011011110111001010101110000010111000); #20
	MCMC_indirect_write(11'd704, 68'b01011000000000000010110000000000000101100000000000001011000000000000); #20
	MCMC_indirect_write(11'd705, 68'b01001110101001100010100101110011000101110000010111101010111001100101); #20
	MCMC_indirect_write(11'd706, 68'b01011001001110001010000100100010000100010001111010101001000111111110); #20
	MCMC_indirect_write(11'd707, 68'b01100110011011111011000111010110000100000100011100101101110111001101); #20
	MCMC_indirect_write(11'd708, 68'b00101101111100000011000100100001010110000011100111101110110011011111); #20
	MCMC_indirect_write(11'd709, 68'b10000101000010110011110001101001100101001000010000001011011011001011); #20
	MCMC_indirect_write(11'd710, 68'b00000001000010100000001110000111010010101001111010100101110001110100); #20
	MCMC_indirect_write(11'd711, 68'b01011101101111111010111100010111110110000000010001001011011011111100); #20
	MCMC_indirect_write(11'd712, 68'b10001101011101100101001001101110011100010111000010111000011101000001); #20
	MCMC_indirect_write(11'd713, 68'b01001100000001010011010110110000110100111110001100001110111011111001); #20
	MCMC_indirect_write(11'd714, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd715, 68'b10010111101010110100100001100110101001001100001000101101001110010001); #20
	MCMC_indirect_write(11'd716, 68'b10110110110100101100011101010010101001110100000100001110001100110011); #20
	MCMC_indirect_write(11'd717, 68'b00010100110110010000000000000000000001110101011100100011001111110000); #20
	MCMC_indirect_write(11'd718, 68'b01010001000111111010000001101011000101110000110101001010011111011111); #20
	MCMC_indirect_write(11'd719, 68'b01000001101101100001110111111000100011010111001110001011000100011001); #20
	MCMC_indirect_write(11'd720, 68'b10101000110001100110010011001110011111000010111111111110010110010001); #20
	MCMC_indirect_write(11'd721, 68'b01000001010011100001011001010101100001110011000101000111111011001001); #20
	MCMC_indirect_write(11'd722, 68'b00000110100010000000000000000000000001100011111101000000000000000000); #20
	MCMC_indirect_write(11'd723, 68'b01010001011100010011000011100101000110001001001010001001010110011001); #20
	MCMC_indirect_write(11'd724, 68'b00100011011100000000111110101101010001101001000011100100010000101111); #20
	MCMC_indirect_write(11'd725, 68'b10010011111111010100010000110001010101111101111000100111111000001011); #20
	MCMC_indirect_write(11'd726, 68'b10000000110110001011100000001000010110110111100100001100010000110101); #20
	MCMC_indirect_write(11'd727, 68'b10000011111000100011110001011100100110011010110110100110111011010011); #20
	MCMC_indirect_write(11'd728, 68'b00001000010111101000000000000000000000011100111001000010011101000011); #20
	MCMC_indirect_write(11'd729, 68'b01111110000100010100001100110011000111011000001011001011011000100001); #20
	MCMC_indirect_write(11'd730, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd731, 68'b00000000000000000000000000000000000000000000000000000001011101110101); #20
	MCMC_indirect_write(11'd732, 68'b11111110111110110111110110011110101110010101100101111111010101001010); #20
	MCMC_indirect_write(11'd733, 68'b01000101111110110011000100011101011000111001110000010000101101101000); #20
	MCMC_indirect_write(11'd734, 68'b11011000011000101110100100111101101101000111100001111011000001110110); #20
	MCMC_indirect_write(11'd735, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd736, 68'b00111001111011111001111011001100100010111101111011001001000101011010); #20
	MCMC_indirect_write(11'd737, 68'b01010111000100100010010100100101000010101000100001000101000101001101); #20
	MCMC_indirect_write(11'd738, 68'b00100001000001010010101011111000010101100111000100110010110000010000); #20
	MCMC_indirect_write(11'd739, 68'b01000001101100001010110010001011100111101010000101101100100100011111); #20
	MCMC_indirect_write(11'd740, 68'b11000000100001111100101101011100111011011001010011001111110101000111); #20
	MCMC_indirect_write(11'd741, 68'b00001010000101000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd742, 68'b01110101111010011011010010110010110110000010101101101011000101011011); #20
	MCMC_indirect_write(11'd743, 68'b00000000000000000000000000000000000000000010001011000001011011111101); #20
	MCMC_indirect_write(11'd744, 68'b11111110101100000111001000000100001101100010100100011100110100001100); #20
	MCMC_indirect_write(11'd745, 68'b01100011101101010010101100000011110110110100000101001111011111010011); #20
	MCMC_indirect_write(11'd746, 68'b00000000000000000000000000000000000010001100101010000000111101111111); #20
	MCMC_indirect_write(11'd747, 68'b10000100100100111100100110010100011001010101010000010000011111011000); #20
	MCMC_indirect_write(11'd748, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd749, 68'b01011111100001110010001001001101110100011010111011000111011001001100); #20
	MCMC_indirect_write(11'd750, 68'b10111011010011101110010101010101101011001000011000011000010111111001); #20
	MCMC_indirect_write(11'd751, 68'b00110010011011111010110010001100010100110111011010100111010001110010); #20
	MCMC_indirect_write(11'd752, 68'b01010100000000000010111101101111010111000001101001101111111101101000); #20
	MCMC_indirect_write(11'd753, 68'b00001100000110010001100101101001010011010111100110100111011010001000); #20
	MCMC_indirect_write(11'd754, 68'b11101111010101001101111000011100001100011000000111111000110011001110); #20
	MCMC_indirect_write(11'd755, 68'b01100101001011010011101010001001000111100111100100110001001101010010); #20
	MCMC_indirect_write(11'd756, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd757, 68'b01000001110010100010111101111101110101100110010100000101111001110011); #20
	MCMC_indirect_write(11'd758, 68'b01000110010100110011010101010101100101001101011010001010000010001011); #20
	MCMC_indirect_write(11'd759, 68'b10000100100111111100101001010010001001101001100001110110111110110100); #20
	MCMC_indirect_write(11'd760, 68'b00111101000100110001111111010010010011100110001100000100111100101111); #20
	MCMC_indirect_write(11'd761, 68'b01001100100000011001110001010011100010010101111110100100010111110010); #20
	MCMC_indirect_write(11'd762, 68'b01111111110100011011001010101110100111011010011110010000111100101010); #20
	MCMC_indirect_write(11'd763, 68'b01011101000100011001111011001100110010010100001110000100100000100101); #20
	MCMC_indirect_write(11'd764, 68'b01001111101010001001000000011100010000000000000000000001111010111101); #20
	MCMC_indirect_write(11'd765, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd766, 68'b00011100110111101000101010110101110001001101111001100011100110110001); #20
	MCMC_indirect_write(11'd767, 68'b10100011000000000101000001010010101000101001010100110001111111000110); #20
	MCMC_indirect_write(11'd768, 68'b01100000000000000011000000000000000110000000000000001100000000000000); #20
	MCMC_indirect_write(11'd769, 68'b01011111100101100010110100001010000101101100111001101100110110000101); #20
	MCMC_indirect_write(11'd770, 68'b01100101001111010011100001111010000101001110100010101010111011100000); #20
	MCMC_indirect_write(11'd771, 68'b10001111010110000011111011111100001000001000001110101011110111001000); #20
	MCMC_indirect_write(11'd772, 68'b01111110010011110011001100110000100101010001011001001100010111011001); #20
	MCMC_indirect_write(11'd773, 68'b10010010000111000011101011001111110011010111010111000011001011100000); #20
	MCMC_indirect_write(11'd774, 68'b10110010100001011100111101111000101010000111101111110011000010010010); #20
	MCMC_indirect_write(11'd775, 68'b01011111011101000011111101001011011001011101110110010011110011100010); #20
	MCMC_indirect_write(11'd776, 68'b00010111110001010001000100010100010011000010101000100011001111101000); #20
	MCMC_indirect_write(11'd777, 68'b00100001111011111000101011000001000101001000110010101011100011000001); #20
	MCMC_indirect_write(11'd778, 68'b01010100110000110010111101101000110100001111011110000111101001010001); #20
	MCMC_indirect_write(11'd779, 68'b10101011100100110110010101100000101111000111000100111011011101000110); #20
	MCMC_indirect_write(11'd780, 68'b00000000000000000000000000000000000000111101101101100000000000000000); #20
	MCMC_indirect_write(11'd781, 68'b00000000000000000000000000000000000000001000010011000000000000000000); #20
	MCMC_indirect_write(11'd782, 68'b10000101010001100011101100100111010111111010011100001110000001101001); #20
	MCMC_indirect_write(11'd783, 68'b01011111100010111100100011110110001010010100000000111010011011110111); #20
	MCMC_indirect_write(11'd784, 68'b01110010011001001011101101111011101000000100101110010001011011011011); #20
	MCMC_indirect_write(11'd785, 68'b01110101100010101011011110011111100111100010100111101011111101001000); #20
	MCMC_indirect_write(11'd786, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd787, 68'b10010111101110011101010001000010011010011100101100011000000001101011); #20
	MCMC_indirect_write(11'd788, 68'b10011000000001010011101000101010100110110111011100110101011101010011); #20
	MCMC_indirect_write(11'd789, 68'b01111101101111000011100110000010010110010111111100101110100000111001); #20
	MCMC_indirect_write(11'd790, 68'b00111010100001101000111000010010100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd791, 68'b10101101010001001101110001000001111010010001110000111011000110111001); #20
	MCMC_indirect_write(11'd792, 68'b01101000000001000010011010000110010110010110000010101111010010000010); #20
	MCMC_indirect_write(11'd793, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd794, 68'b01011001001001000010101101101100000110110001001100001101011000111001); #20
	MCMC_indirect_write(11'd795, 68'b01110100111000001011111111000110011000000100100111110000110101011101); #20
	MCMC_indirect_write(11'd796, 68'b00000111010101000000000000000000000001010111101111100000011001000110); #20
	MCMC_indirect_write(11'd797, 68'b00111010110101010010001110111001010110101001000110001011110011100111); #20
	MCMC_indirect_write(11'd798, 68'b10000000000000000010000000000000000111100010001101010000000000000000); #20
	MCMC_indirect_write(11'd799, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd800, 68'b10101010100101001101000111011010100111101001101100001011100000011001); #20
	MCMC_indirect_write(11'd801, 68'b01010101000111011011001010000001100110101111001010101111110010001011); #20
	MCMC_indirect_write(11'd802, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd803, 68'b00000100010101100000110010110111110011001101001100100111100110101110); #20
	MCMC_indirect_write(11'd804, 68'b01101110001101010011101111110011010101000001001001001101001100001000); #20
	MCMC_indirect_write(11'd805, 68'b10001011010110010011101001101001000101101011001111001101101001011101); #20
	MCMC_indirect_write(11'd806, 68'b10000000000000000100000000000000001111011011011101111010011101111000); #20
	MCMC_indirect_write(11'd807, 68'b00000000000000000000000000000000000000001011110011100010110000111001); #20
	MCMC_indirect_write(11'd808, 68'b01000011001000110010011011010011110111010111100101101011110110100101); #20
	MCMC_indirect_write(11'd809, 68'b11001011010011100111011000010110001111100001001110011100101110010110); #20
	MCMC_indirect_write(11'd810, 68'b10010111000110010101001000110101011000101101101111101111001100111110); #20
	MCMC_indirect_write(11'd811, 68'b00111100010111110001010110111011110101001001100100101011101011110010); #20
	MCMC_indirect_write(11'd812, 68'b00111000000000101001010100000101100000100001010011000100000110010100); #20
	MCMC_indirect_write(11'd813, 68'b10000000110111001011111100111111011001000001100110010011100011000000); #20
	MCMC_indirect_write(11'd814, 68'b00100110010000000001111010001101110011011000011100100100000101001111); #20
	MCMC_indirect_write(11'd815, 68'b01110100111011111100001100100001110110111000111101101110010001110000); #20
	MCMC_indirect_write(11'd816, 68'b01100010011110111101001011111011101100001011100110011010001101000101); #20
	MCMC_indirect_write(11'd817, 68'b00111000100111110010011000001100110011100000110111001000110001111101); #20
	MCMC_indirect_write(11'd818, 68'b00110001101100100001110001011001000010100001100110100100110110000011); #20
	MCMC_indirect_write(11'd819, 68'b11100110001010110110111010110011111011101011001010111101000101110000); #20
	MCMC_indirect_write(11'd820, 68'b11000111100000010101100010111111011001110011100001010100000110000000); #20
	MCMC_indirect_write(11'd821, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd822, 68'b00010111100000010001011111100101110010000000000100000010100010001101); #20
	MCMC_indirect_write(11'd823, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd824, 68'b01111101000100000100010110100001100111010111110111101111000110111000); #20
	MCMC_indirect_write(11'd825, 68'b00111011011100111001011101000000010011101110011111101000101001001110); #20
	MCMC_indirect_write(11'd826, 68'b00110011110001001001111001010110000101010101111010101011110011011001); #20
	MCMC_indirect_write(11'd827, 68'b00110011100100011001101111000110010010100100111010101000101000111110); #20
	MCMC_indirect_write(11'd828, 68'b10010111101000101100010101100100101000011100101111101010110110100111); #20
	MCMC_indirect_write(11'd829, 68'b10000001010011100100011100010011001000111000110100010010010100101111); #20
	MCMC_indirect_write(11'd830, 68'b01001101111110001010001011000001100011110101111001100100001001010011); #20
	MCMC_indirect_write(11'd831, 68'b01001110100010000011000000011100000101001000100100001100001110100001); #20
	MCMC_indirect_write(11'd832, 68'b01101000000000000011010000000000000110100000000000001101000000000000); #20
	MCMC_indirect_write(11'd833, 68'b01101010010110111011001101011011000110011100100110001011111100101110); #20
	MCMC_indirect_write(11'd834, 68'b01101001010011011011000011111110010110110110110110101111010110010001); #20
	MCMC_indirect_write(11'd835, 68'b01110111000010110011000111001111110111111011010000001101111011100011); #20
	MCMC_indirect_write(11'd836, 68'b01011001011001000010110110011001100101100110011000001101111010011110); #20
	MCMC_indirect_write(11'd837, 68'b01011101100110111011101110000101101000001110111000010100001001111100); #20
	MCMC_indirect_write(11'd838, 68'b00101000101000110010101101111011100001001111000000000001011001001100); #20
	MCMC_indirect_write(11'd839, 68'b10000010001000000011110111011101100110001011000011100110111001111101); #20
	MCMC_indirect_write(11'd840, 68'b10111001010100001101111010110100011101010010110110111010010011010000); #20
	MCMC_indirect_write(11'd841, 68'b01000001111110100011000001101011110101100111101001001100111000000000); #20
	MCMC_indirect_write(11'd842, 68'b00110000111010101010000010000001010011100110100100000110100001010110); #20
	MCMC_indirect_write(11'd843, 68'b00100010101011000001100001100100000100000001000000101000010010111000); #20
	MCMC_indirect_write(11'd844, 68'b11010110011111111101110010111101011101000000011010010110101000011110); #20
	MCMC_indirect_write(11'd845, 68'b10000000000000000011101011000010111111000111010000111011101101000001); #20
	MCMC_indirect_write(11'd846, 68'b01000110100010001010010000101011110010001001000100000110001101000111); #20
	MCMC_indirect_write(11'd847, 68'b01001111100111111011011010001010001000110001001000110100000011011010); #20
	MCMC_indirect_write(11'd848, 68'b01101101111000100100010100101100111001000011110110010010000001100001); #20
	MCMC_indirect_write(11'd849, 68'b10010101111011001011000100001110000100101101110100100111000011001111); #20
	MCMC_indirect_write(11'd850, 68'b11011000010100111111100011110101011110011000001100111011010011000010); #20
	MCMC_indirect_write(11'd851, 68'b00000000000000000000100000110010100011101010100101000000111111100001); #20
	MCMC_indirect_write(11'd852, 68'b00101010100110000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd853, 68'b01001000111100101010000010111011010100110001010100100100001100011011); #20
	MCMC_indirect_write(11'd854, 68'b10011110110010010101000010001111000111111111111101001100110101101010); #20
	MCMC_indirect_write(11'd855, 68'b10111001110011010100100111101101001000100110100100110100111100000101); #20
	MCMC_indirect_write(11'd856, 68'b00110011001111001001011001000000110011101101111111100011001111111010); #20
	MCMC_indirect_write(11'd857, 68'b01101100001101001100000010011000000111101100011001001100011101010001); #20
	MCMC_indirect_write(11'd858, 68'b10100100110011000011010011100011110111111111010110001110001110011001); #20
	MCMC_indirect_write(11'd859, 68'b01000101011001000010101100100111010101010100111100001001111101000000); #20
	MCMC_indirect_write(11'd860, 68'b01111010111101011101101010111100111011010000111111110101011111001111); #20
	MCMC_indirect_write(11'd861, 68'b10011001111110100011101110111110000111110101111110101101001110011010); #20
	MCMC_indirect_write(11'd862, 68'b11000010000000001110010110011110011111000001011101011110011001111000); #20
	MCMC_indirect_write(11'd863, 68'b01110010110000101000111110010100010011000011000110100101100001111101); #20
	MCMC_indirect_write(11'd864, 68'b11011100001010101110101101011101111100000100100110110111000100111110); #20
	MCMC_indirect_write(11'd865, 68'b01101010100100111011101101011100000100101110101101101110001110111111); #20
	MCMC_indirect_write(11'd866, 68'b01100101010001010011110010111000111000010011101010101111110001011111); #20
	MCMC_indirect_write(11'd867, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd868, 68'b00111000001110100001100111110010110010101101011001100111011001101101); #20
	MCMC_indirect_write(11'd869, 68'b01001000101101110011000001001011100111001000111000001110011110111001); #20
	MCMC_indirect_write(11'd870, 68'b10011000001001100100110100110010011001110010010100010011001100001110); #20
	MCMC_indirect_write(11'd871, 68'b10001110101110001100110100101110011001001110000010010001000100101101); #20
	MCMC_indirect_write(11'd872, 68'b10111010100101110110000111001100001101101101110101111000000011000111); #20
	MCMC_indirect_write(11'd873, 68'b11010001111101100110001100001101011010101000011010111101011100111010); #20
	MCMC_indirect_write(11'd874, 68'b01010000011000111001110000001011100010010010010101100010100110110100); #20
	MCMC_indirect_write(11'd875, 68'b10000000000000001000000000000000010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd876, 68'b00100001001001110000111100001001110010100110000111100101001100000001); #20
	MCMC_indirect_write(11'd877, 68'b01000101010111111010101000010000000010110111001001100011011011011110); #20
	MCMC_indirect_write(11'd878, 68'b10011010001000101011000000011001100110000100010001001111010001110110); #20
	MCMC_indirect_write(11'd879, 68'b00111111110101110011000001101011110101011100100010101101101101011011); #20
	MCMC_indirect_write(11'd880, 68'b01010111110101000011000000110101110011111101010110001011001001111101); #20
	MCMC_indirect_write(11'd881, 68'b10000000000000000100000000000000001111010101010101100000000000000000); #20
	MCMC_indirect_write(11'd882, 68'b10010010100111000101101011000100111011011110111000010000000001101001); #20
	MCMC_indirect_write(11'd883, 68'b01101110010110011100001110100011111001001010111111110000111101011101); #20
	MCMC_indirect_write(11'd884, 68'b00101110101011011001110100101110010010111011101000100111111010100110); #20
	MCMC_indirect_write(11'd885, 68'b11001001011100111101111011100110001001110001100110010101100001110101); #20
	MCMC_indirect_write(11'd886, 68'b10010111100101110011011100110100100110101010011100101111000110001000); #20
	MCMC_indirect_write(11'd887, 68'b10110100011000100110010010011101101100110111000010011011111101000001); #20
	MCMC_indirect_write(11'd888, 68'b11000011111100101110100000100100001101100111110010110111100100001101); #20
	MCMC_indirect_write(11'd889, 68'b01111011010100110100110110100011001000011011011111010010101100000111); #20
	MCMC_indirect_write(11'd890, 68'b10001101110111011100110001111010101010000011101111010100110110001111); #20
	MCMC_indirect_write(11'd891, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd892, 68'b01010011010001101011001110000101000101111001010101001001111011011111); #20
	MCMC_indirect_write(11'd893, 68'b10101110111110101011110000111100011001111011010101010100010111101011); #20
	MCMC_indirect_write(11'd894, 68'b01100110111110000011101111010111010111111110001000110001010100011110); #20
	MCMC_indirect_write(11'd895, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd896, 68'b01110000000000000011100000000000000111000000000000001110000000000000); #20
	MCMC_indirect_write(11'd897, 68'b01111000001001110011010111000111110110011100100000001100000111100110); #20
	MCMC_indirect_write(11'd898, 68'b01011011100001101010101011111000100110111010100011001011111001101000); #20
	MCMC_indirect_write(11'd899, 68'b10011100011001100011110110110000100110100111100001001011000100101001); #20
	MCMC_indirect_write(11'd900, 68'b01101110000101111011001011100000010111101100000011001011101010101000); #20
	MCMC_indirect_write(11'd901, 68'b01011110111000110011010010101001101000100011011101010011000001011101); #20
	MCMC_indirect_write(11'd902, 68'b10000001111010001011110111100101011000110101110100110001000001101110); #20
	MCMC_indirect_write(11'd903, 68'b11000000100101010100001001110111011000100110011011110001111100101101); #20
	MCMC_indirect_write(11'd904, 68'b10000000000000000111101110111111001000000000000000011110010011011100); #20
	MCMC_indirect_write(11'd905, 68'b10101010111100100101010000000011011001000100011000101111001110000110); #20
	MCMC_indirect_write(11'd906, 68'b11011111100000011110111101001011110000000000000000011100101101000011); #20
	MCMC_indirect_write(11'd907, 68'b01100010001011000010100000110110100101100001101010001101011001111110); #20
	MCMC_indirect_write(11'd908, 68'b01110100101001000100101000001110011000100101010101001101000101110100); #20
	MCMC_indirect_write(11'd909, 68'b10001011000111101010101100000000010011011101011011100111101100100010); #20
	MCMC_indirect_write(11'd910, 68'b10001100000011011011010100111011000110001100110100101101110011110010); #20
	MCMC_indirect_write(11'd911, 68'b00101000001110011000110000011010010010011001101101000011110100010001); #20
	MCMC_indirect_write(11'd912, 68'b01100011000010101011011011111000101000000011101111010110000011001011); #20
	MCMC_indirect_write(11'd913, 68'b01100001111101100011010010100000110101101010011001101010111110110111); #20
	MCMC_indirect_write(11'd914, 68'b11110110011110101000000000000000001111101010111100011110110000101111); #20
	MCMC_indirect_write(11'd915, 68'b10111000010110011110001110011001111011100000100101111010110100110110); #20
	MCMC_indirect_write(11'd916, 68'b00101100001110011010010001000101110011100011111111101001000111100111); #20
	MCMC_indirect_write(11'd917, 68'b00101001011010100000111101011000100001001110110110100000000000000000); #20
	MCMC_indirect_write(11'd918, 68'b01001000101010111010011101000010110101111111000111001100001011101110); #20
	MCMC_indirect_write(11'd919, 68'b11001110100101001100001001011010011101101110010001100000000000000000); #20
	MCMC_indirect_write(11'd920, 68'b10000111110101010010010111011110110001101011010101100001110100110111); #20
	MCMC_indirect_write(11'd921, 68'b00110011011111111001100011000011010101000000111100000111001001111111); #20
	MCMC_indirect_write(11'd922, 68'b01000011010101011001000101010011110011110011011000100111100110111011); #20
	MCMC_indirect_write(11'd923, 68'b11011011110010110101101100101101001001000011101000110101010100100001); #20
	MCMC_indirect_write(11'd924, 68'b11110010111110110000000000000000010000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd925, 68'b00100101001111011010010101100010000110010000000010010001000010111101); #20
	MCMC_indirect_write(11'd926, 68'b10010100101001010101011111100001011010111100100100011001110000010010); #20
	MCMC_indirect_write(11'd927, 68'b10011011011010001100101000010101011010110100100011110110111000101010); #20
	MCMC_indirect_write(11'd928, 68'b01000101110111010010111010111010000101011011110110001001100010010111); #20
	MCMC_indirect_write(11'd929, 68'b01101000110111001100110110100100110111101001110100110000001101110000); #20
	MCMC_indirect_write(11'd930, 68'b01101100011101111100010101111010101000111010100011101110001011100101); #20
	MCMC_indirect_write(11'd931, 68'b01100001001110100010110111110000010101001111000111101111110111010001); #20
	MCMC_indirect_write(11'd932, 68'b10100001111001011111010010111000011101110011101111111001110101001010); #20
	MCMC_indirect_write(11'd933, 68'b10110001110010111110100010010111111101001011001111011100010101100000); #20
	MCMC_indirect_write(11'd934, 68'b11010101111011000111100001101000110000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd935, 68'b01011001000101101001110001011110000001101101000011100000000000000000); #20
	MCMC_indirect_write(11'd936, 68'b00001011100000111000000000000000000001000101110101100011111011011100); #20
	MCMC_indirect_write(11'd937, 68'b00000000000000000000101010110111100000110110011010100101110011101010); #20
	MCMC_indirect_write(11'd938, 68'b00111100010101000001111010001110110101001101110000100100101010110001); #20
	MCMC_indirect_write(11'd939, 68'b11010101011011001101111101101111001010110111001000110100111100000110); #20
	MCMC_indirect_write(11'd940, 68'b10011011000011010101001111100010011100110110000011011001101111010100); #20
	MCMC_indirect_write(11'd941, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd942, 68'b01010011100000001010100011110111110101101110111101101010000111111001); #20
	MCMC_indirect_write(11'd943, 68'b00110100001101001000101101111001100001010000011100000000000000000000); #20
	MCMC_indirect_write(11'd944, 68'b10100001101011010110101101011111010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd945, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd946, 68'b10100010101101101100111110010011111101101011101011111000111110010011); #20
	MCMC_indirect_write(11'd947, 68'b10100001001110001110001010110000001110010111110101111011101100000001); #20
	MCMC_indirect_write(11'd948, 68'b10100111100010101110011111101100101011111000011110111001001101010011); #20
	MCMC_indirect_write(11'd949, 68'b10101110111010001100101011111110110111010000001001101101000000110010); #20
	MCMC_indirect_write(11'd950, 68'b10101011100011101101011110011000111000000111000000110100001001101000); #20
	MCMC_indirect_write(11'd951, 68'b11001100011110001101110100011110011100000101110101111100010111100111); #20
	MCMC_indirect_write(11'd952, 68'b01000000011001011010010001111111110101110101110101100111101001010111); #20
	MCMC_indirect_write(11'd953, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd954, 68'b01111110001111010101101011010001111011101110100010111011001000110000); #20
	MCMC_indirect_write(11'd955, 68'b01110100001111100011111001011001100111101011011000101111101010101100); #20
	MCMC_indirect_write(11'd956, 68'b11000111000111111110011011000011101101101000111010010110011111001011); #20
	MCMC_indirect_write(11'd957, 68'b01010111110000100011101011110000111010100000110111111000010110010111); #20
	MCMC_indirect_write(11'd958, 68'b01110001000111010010100000110010000101011111111111101110001001100000); #20
	MCMC_indirect_write(11'd959, 68'b01111001110101110100110010110010110111010011001110001111111010110011); #20
	MCMC_indirect_write(11'd960, 68'b01111000000000000011110000000000000111100000000000001111000000000000); #20
	MCMC_indirect_write(11'd961, 68'b01111111001001011100000001101001110111101101100010101110100101010101); #20
	MCMC_indirect_write(11'd962, 68'b01110101100000100011101000100000000111101000111010001100110001111001); #20
	MCMC_indirect_write(11'd963, 68'b10000100011010111100001101111011011000100010010100101011100001011010); #20
	MCMC_indirect_write(11'd964, 68'b01100100111101011100010100100101000111111010010010110000010000001111); #20
	MCMC_indirect_write(11'd965, 68'b00111111111001100010110010111101110111110111100110010000101100000111); #20
	MCMC_indirect_write(11'd966, 68'b01011100101110010011000101111101010110001111011001101011110001111101); #20
	MCMC_indirect_write(11'd967, 68'b01110101001011010101100010110110011010011100010101010110010110011101); #20
	MCMC_indirect_write(11'd968, 68'b10100000101100000101110010110001101100100011101001010101011000010101); #20
	MCMC_indirect_write(11'd969, 68'b10001000111011100101010100100111011010101110010101011100000001001010); #20
	MCMC_indirect_write(11'd970, 68'b01101011001011111011110000010110010111100011110011001011010101001000); #20
	MCMC_indirect_write(11'd971, 68'b10111010010000010110011001101100111011001001110101010100000111010100); #20
	MCMC_indirect_write(11'd972, 68'b01110000001100100100000010011001110111110100011111010011010100111101); #20
	MCMC_indirect_write(11'd973, 68'b10100000100000101011101000101011010111010011101100001110100010100110); #20
	MCMC_indirect_write(11'd974, 68'b01000011101011010010110000000111000111110001111100001101000000000111); #20
	MCMC_indirect_write(11'd975, 68'b01011100111100100010001101111010110100110011101100001100000110110001); #20
	MCMC_indirect_write(11'd976, 68'b01111101101100100110000100001011001100110100101010111001111111001000); #20
	MCMC_indirect_write(11'd977, 68'b10101001100111011011101110111111000101110110001111110000101011000001); #20
	MCMC_indirect_write(11'd978, 68'b01111000110101111100111101001001001001101101100101010111001011100010); #20
	MCMC_indirect_write(11'd979, 68'b10001001101001111100100111011010011010010010111001110101000000011110); #20
	MCMC_indirect_write(11'd980, 68'b00100100110001011000111001011000010011000110111011100000000000000000); #20
	MCMC_indirect_write(11'd981, 68'b01101111000000010100101010111010111010001010111111110100001000001110); #20
	MCMC_indirect_write(11'd982, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd983, 68'b01001011110010111001110110110001010001111110001111000010110001100010); #20
	MCMC_indirect_write(11'd984, 68'b10010011101110010100011011101100111001011010011001101110010111011101); #20
	MCMC_indirect_write(11'd985, 68'b10110110001000010111001000111011101110101110110000011111011001111010); #20
	MCMC_indirect_write(11'd986, 68'b01011000100000101011011001110000000101110101011111101100000010101011); #20
	MCMC_indirect_write(11'd987, 68'b10100000111010100101011000111000001010110001111101010011101011011100); #20
	MCMC_indirect_write(11'd988, 68'b01000001000000110001110100110000010000111011010110100000100111101110); #20
	MCMC_indirect_write(11'd989, 68'b10010111100101011100001010110011001011001100011100011101110011101101); #20
	MCMC_indirect_write(11'd990, 68'b01111111000000110011100101010111100111010111111010001110011101010111); #20
	MCMC_indirect_write(11'd991, 68'b01001000010111001001010101000001010000100111011100100011010000001001); #20
	MCMC_indirect_write(11'd992, 68'b10011110111010111010110100100001000101110000110101001000010111101110); #20
	MCMC_indirect_write(11'd993, 68'b00110010110000101010011001101010110110110001011001101011000011101001); #20
	MCMC_indirect_write(11'd994, 68'b10000010010111101011111101100010001001111101010001110001110111000000); #20
	MCMC_indirect_write(11'd995, 68'b10011010000111111100101101011100010110000101000110001000111111111001); #20
	MCMC_indirect_write(11'd996, 68'b10110010010011111110010001011011111010100010000010011001100001111101); #20
	MCMC_indirect_write(11'd997, 68'b00000110111011011000000000000000000011100010001100000011010100000111); #20
	MCMC_indirect_write(11'd998, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd999, 68'b10101100100110111101010011011110111011001100111011110000100000110011); #20
	MCMC_indirect_write(11'd1000, 68'b10101101010011111100110111010001010101010001110101100100011101111000); #20
	MCMC_indirect_write(11'd1001, 68'b01011001101001110010011000100010001111111111110011100011111110000110); #20
	MCMC_indirect_write(11'd1002, 68'b00001111000100010000011001001001100000000000000000000010100110111000); #20
	MCMC_indirect_write(11'd1003, 68'b10000110010010010100100010101000000111010111111011000011100110101010); #20
	MCMC_indirect_write(11'd1004, 68'b11110100100100100100000000000000011011001010111111110011110001010100); #20
	MCMC_indirect_write(11'd1005, 68'b11010001010101111110000111101010011111001000010110111010000110011110); #20
	MCMC_indirect_write(11'd1006, 68'b01010101001000100001110110010001110011110011111100000011010010000010); #20
	MCMC_indirect_write(11'd1007, 68'b01011001010111011001110001010100100011010101000001010001000111100100); #20
	MCMC_indirect_write(11'd1008, 68'b10000000000000001111000010011111100000000000000001000000000000000000); #20
	MCMC_indirect_write(11'd1009, 68'b10001100001110010111111010010001001110111111100011011010110000010100); #20
	MCMC_indirect_write(11'd1010, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1011, 68'b01110000101111100111001000001000101101110000100111010001011001001110); #20
	MCMC_indirect_write(11'd1012, 68'b10101011010010110100100010000111010101010000111111101100100001101100); #20
	MCMC_indirect_write(11'd1013, 68'b10101001110111010100010001000111100111001100011100010101001001010000); #20
	MCMC_indirect_write(11'd1014, 68'b10000101000011100010111100111000110101110011001101001000111000011110); #20
	MCMC_indirect_write(11'd1015, 68'b10001001011101011100000001110010110110010101011101101101011101100100); #20
	MCMC_indirect_write(11'd1016, 68'b00000000000000000000001011000010110000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1017, 68'b11100011011101001111010011101010111110010011010001110010010111101100); #20
	MCMC_indirect_write(11'd1018, 68'b01001111110011010101010000101111001000000011111010001101111011100110); #20
	MCMC_indirect_write(11'd1019, 68'b00111111111000111011000001111101110101001000010000100111110011100110); #20
	MCMC_indirect_write(11'd1020, 68'b11010111101011011111110110001001010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1021, 68'b00011100000110100001000001101110000010111100111110100110100011110110); #20
	MCMC_indirect_write(11'd1022, 68'b01111100111001111100011001001010001011100000100001011001001010011000); #20
	MCMC_indirect_write(11'd1023, 68'b01100001100000001010000001011101010011010110100100001100100011111110); #20
	MCMC_indirect_write(11'd1024, 68'b10000000000000000100000000000000001000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1025, 68'b10000000000001010011101110111101000111111011010101011100001010100000); #20
	MCMC_indirect_write(11'd1026, 68'b10000011011011111000101100000110010000110110100001011111111100110100); #20
	MCMC_indirect_write(11'd1027, 68'b01110100110001100011101100110010000101101110110010101111100011101010); #20
	MCMC_indirect_write(11'd1028, 68'b10001101110010000100100011000010011010000000101001110110101001110010); #20
	MCMC_indirect_write(11'd1029, 68'b10001010010011110101011110010011011001100110111011011101010010101010); #20
	MCMC_indirect_write(11'd1030, 68'b10010001001000010100010010011000001111001101111101100001100111010110); #20
	MCMC_indirect_write(11'd1031, 68'b10000101011000000101010000001110010111111000000100100110010000100100); #20
	MCMC_indirect_write(11'd1032, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1033, 68'b10111111100010101011010001101111011011000110101010110101101011011100); #20
	MCMC_indirect_write(11'd1034, 68'b01101111111110111011100100100001010110111110001010110111011101010000); #20
	MCMC_indirect_write(11'd1035, 68'b01001100011010101011001011101000010110110001000111100010001110010000); #20
	MCMC_indirect_write(11'd1036, 68'b11001101111100101110010101100111001010100100111110100010100110011110); #20
	MCMC_indirect_write(11'd1037, 68'b10000000000000000100000000000000011111110101000011111100111011010000); #20
	MCMC_indirect_write(11'd1038, 68'b10101101001000001101100011010110111011011100000100101100101101101100); #20
	MCMC_indirect_write(11'd1039, 68'b01011110001101000100010011111111011000011001111100101111110010001110); #20
	MCMC_indirect_write(11'd1040, 68'b10001001001111011011000101011101010110011010011100101010001001011100); #20
	MCMC_indirect_write(11'd1041, 68'b01000010011100001010000110000101100101111110111110011010010100100010); #20
	MCMC_indirect_write(11'd1042, 68'b10001011010111010100011110010011010110010101101100100001101001100000); #20
	MCMC_indirect_write(11'd1043, 68'b00011000101100111001100001010100000001110001110111100011100100011000); #20
	MCMC_indirect_write(11'd1044, 68'b10000111100100111101010000110001011000100111000111101101001010010000); #20
	MCMC_indirect_write(11'd1045, 68'b10100110110101001011101000100110011001110111110001101101111010111000); #20
	MCMC_indirect_write(11'd1046, 68'b01110011000001100101110110000011000111111010011011010001001100110010); #20
	MCMC_indirect_write(11'd1047, 68'b10101111100100010101011001110001101001001101001100100111100111100100); #20
	MCMC_indirect_write(11'd1048, 68'b01100010100001001010100101101111010100011001111000101011100010000010); #20
	MCMC_indirect_write(11'd1049, 68'b01110011010001111100100101010000011010110010111110101101000011111010); #20
	MCMC_indirect_write(11'd1050, 68'b10011011100111101001111100111010010000111001000011011111101100000110); #20
	MCMC_indirect_write(11'd1051, 68'b11101000000101010110011001000100101010000111111100110011110110000000); #20
	MCMC_indirect_write(11'd1052, 68'b10001011100000110100100011001010110111010001010110011111110011011110); #20
	MCMC_indirect_write(11'd1053, 68'b10101111110101001110010011100101101101101001001110110000011100010100); #20
	MCMC_indirect_write(11'd1054, 68'b11010100011100111111010100100100011100011011000110101100101011110100); #20
	MCMC_indirect_write(11'd1055, 68'b10110011000010001101110001011001111000000111010001100111000011010100); #20
	MCMC_indirect_write(11'd1056, 68'b11010000000101001101111001010111111010101111000001100110110111110110); #20
	MCMC_indirect_write(11'd1057, 68'b00111001001100001011001010000000000100100010010000001110011010100000); #20
	MCMC_indirect_write(11'd1058, 68'b10001010111100011100100000111010010111010001101111010001011000110100); #20
	MCMC_indirect_write(11'd1059, 68'b10010110110111100100101100010111101010000100001101010010111111011000); #20
	MCMC_indirect_write(11'd1060, 68'b11001001100010011110100101111101001110101100010010110001000000000100); #20
	MCMC_indirect_write(11'd1061, 68'b10000001100100100010110001011011001110111110010111100011101000001100); #20
	MCMC_indirect_write(11'd1062, 68'b10101111111111001101011001010101010101111111100110100110000001001100); #20
	MCMC_indirect_write(11'd1063, 68'b10101110000111000101010101111111110110001110110100110010010101111010); #20
	MCMC_indirect_write(11'd1064, 68'b10010100101111001101101111000000111100001100010100100000000000000000); #20
	MCMC_indirect_write(11'd1065, 68'b11101000101001101111111011001000110000000000000000111110011011001110); #20
	MCMC_indirect_write(11'd1066, 68'b01111111010110110111111000100001010000100011010111101010111110110000); #20
	MCMC_indirect_write(11'd1067, 68'b00001100101001000000000000000000000000000000000000000110111001111110); #20
	MCMC_indirect_write(11'd1068, 68'b00110101011010100010110011000010001011110101010011010101011001110010); #20
	MCMC_indirect_write(11'd1069, 68'b01111101110111111101010011001110011010101110001101010111111111110000); #20
	MCMC_indirect_write(11'd1070, 68'b00011111000001101000110100010000000000000011100000100000000000000000); #20
	MCMC_indirect_write(11'd1071, 68'b11110110001000011111101011010000011011101110001100111001010110100100); #20
	MCMC_indirect_write(11'd1072, 68'b10010011111100001011101111011001010110100001000001101001110010001000); #20
	MCMC_indirect_write(11'd1073, 68'b11011111110001101000000000000000010000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1074, 68'b11101001110101011111001100110010101100110000111101101100010100110000); #20
	MCMC_indirect_write(11'd1075, 68'b10000000000000000100000000000000001000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1076, 68'b10000110010110011101010001111100101010001001111000101101000110011000); #20
	MCMC_indirect_write(11'd1077, 68'b10111000010100001110011101010110101100110011101101010100100100100100); #20
	MCMC_indirect_write(11'd1078, 68'b01110010010111100100001111101101001001000010110000110010110111110100); #20
	MCMC_indirect_write(11'd1079, 68'b01001011000101001011100011011000101000000001110010100011011101010110); #20
	MCMC_indirect_write(11'd1080, 68'b10110010000100100101001110010111011010000010011101010000111000010101); #20
	MCMC_indirect_write(11'd1081, 68'b11000110100000010101111011100100001011000100110111010100010101001011); #20
	MCMC_indirect_write(11'd1082, 68'b10000000000000000010000000000000000111100110000000001101100111111011); #20
	MCMC_indirect_write(11'd1083, 68'b10110000101100000100100010100000101100001111010101011010011010101101); #20
	MCMC_indirect_write(11'd1084, 68'b10010110000111001101011000010100001011111110101010010110101011101100); #20
	MCMC_indirect_write(11'd1085, 68'b11101100010001001100000000000000010000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1086, 68'b11100111000000111111111101000101110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1087, 68'b10010000111111100011101000100110001001100110101001110011111110100010); #20
	MCMC_indirect_write(11'd1088, 68'b10001000000000000100010000000000001000100000000000010001000000000000); #20
	MCMC_indirect_write(11'd1089, 68'b01111111000100011011101110111100100111111100101001010010000010011000); #20
	MCMC_indirect_write(11'd1090, 68'b10011101100011100100001010110100101001100010000100010001100110001000); #20
	MCMC_indirect_write(11'd1091, 68'b10000001101011101100010011101100001010010001010011110010011100011001); #20
	MCMC_indirect_write(11'd1092, 68'b01111110000101001011111100010110011001111100100000110010110110011101); #20
	MCMC_indirect_write(11'd1093, 68'b01100101011001011011010101101011101000101011000011110001000000011010); #20
	MCMC_indirect_write(11'd1094, 68'b01100101101101010011010011011010110110001010101001001101101010110111); #20
	MCMC_indirect_write(11'd1095, 68'b10000000000000000011011100000000110111011001110111011110001010001101); #20
	MCMC_indirect_write(11'd1096, 68'b01100111111001001011001110101001000110101010100110101111111111101101); #20
	MCMC_indirect_write(11'd1097, 68'b10011111010010101100111000010111011011111100101110111001111100000011); #20
	MCMC_indirect_write(11'd1098, 68'b10010100001011110101001100000100011101011000011101011000010010111111); #20
	MCMC_indirect_write(11'd1099, 68'b01101011010010011010011100111111000011110101110000001001110001000111); #20
	MCMC_indirect_write(11'd1100, 68'b10101001111101111100100010100000011000000111000101111000101011001101); #20
	MCMC_indirect_write(11'd1101, 68'b01001111101101000010100111111101100111000111100011101110011010101111); #20
	MCMC_indirect_write(11'd1102, 68'b10010011101000100100011101001101110101101101110000101101010001010111); #20
	MCMC_indirect_write(11'd1103, 68'b10111111111001101101001000011000010110111010100000000110101011110111); #20
	MCMC_indirect_write(11'd1104, 68'b10111101011110111110100000000111011101101101100101111010100111101100); #20
	MCMC_indirect_write(11'd1105, 68'b11011110000000101111011001000010101110101011100010011111100101100010); #20
	MCMC_indirect_write(11'd1106, 68'b10010111001011011101010110001111111011110010111100011010111011100100); #20
	MCMC_indirect_write(11'd1107, 68'b01011101110110111010000100110010010001001011111010100110110101110110); #20
	MCMC_indirect_write(11'd1108, 68'b10011010011010001110001011111001011110011000101101011001000001000001); #20
	MCMC_indirect_write(11'd1109, 68'b01000010110111011001110111101100010001101010000101000010000000101010); #20
	MCMC_indirect_write(11'd1110, 68'b10001111101001011010110000110101010101000001110000101001110101101000); #20
	MCMC_indirect_write(11'd1111, 68'b00101000111000011001001101111111100000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1112, 68'b00101111010000111000100110101110000010011001010101000001001111001010); #20
	MCMC_indirect_write(11'd1113, 68'b10011100111000101100001110000000110110000011101100101010010100000010); #20
	MCMC_indirect_write(11'd1114, 68'b01011110000110000010000011100100000011110011011101000110101000101010); #20
	MCMC_indirect_write(11'd1115, 68'b00111100001110010011000001110101010101010101011010101011100011100000); #20
	MCMC_indirect_write(11'd1116, 68'b10110010000000110101001001111010001010000101011100011001011110101110); #20
	MCMC_indirect_write(11'd1117, 68'b01101011100000010011001010011111100111000000110001110001011011101110); #20
	MCMC_indirect_write(11'd1118, 68'b01101111001001101100010101110010011001010000001001110001010111101101); #20
	MCMC_indirect_write(11'd1119, 68'b10011001000110001011110100000111001000010010000101110001011110101001); #20
	MCMC_indirect_write(11'd1120, 68'b11001001011100011111001001001011111111011010111110011011001011111010); #20
	MCMC_indirect_write(11'd1121, 68'b01000000110010110010100011101111100101000010000010001001110000101000); #20
	MCMC_indirect_write(11'd1122, 68'b11100001111111001110110111000010001111100101010010011100101101100100); #20
	MCMC_indirect_write(11'd1123, 68'b10001010000101101101000010010010001010011001101110110111100010101000); #20
	MCMC_indirect_write(11'd1124, 68'b01100000010111000011110111101111011000000101101011001110111111111001); #20
	MCMC_indirect_write(11'd1125, 68'b00000000100111011000000000000000000000000001000010000000101110111100); #20
	MCMC_indirect_write(11'd1126, 68'b10000000111101100100000011100100110101101011010101101110101000001011); #20
	MCMC_indirect_write(11'd1127, 68'b11001101110010000110000010011001011011100010010101011011111010010001); #20
	MCMC_indirect_write(11'd1128, 68'b00110101110111111010111101001011010110100001011001001110110011101101); #20
	MCMC_indirect_write(11'd1129, 68'b10111101010111100101111100100010111101111100011000011001000110000000); #20
	MCMC_indirect_write(11'd1130, 68'b10000000000000000100000000000000001101100111010110011000101111011011); #20
	MCMC_indirect_write(11'd1131, 68'b00000010001100001000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1132, 68'b10010100001100111011000101001001010110010100010010001110100110010110); #20
	MCMC_indirect_write(11'd1133, 68'b11100000001000101110111111111000011011101001010010111010001000111001); #20
	MCMC_indirect_write(11'd1134, 68'b10110101111101100110011011001010111100111110000100111101101110100001); #20
	MCMC_indirect_write(11'd1135, 68'b00100010101100100000001101110111100010010000010011100111110110111110); #20
	MCMC_indirect_write(11'd1136, 68'b11101110111111001111000001110010111111001111100101110000000000000000); #20
	MCMC_indirect_write(11'd1137, 68'b10101101001010100100001011100100010111101110011101010010101101001101); #20
	MCMC_indirect_write(11'd1138, 68'b01110111000111000010101101111001000111010100111100010001011100001101); #20
	MCMC_indirect_write(11'd1139, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1140, 68'b10000101100011011100110000001000001000101001000110110000111011111101); #20
	MCMC_indirect_write(11'd1141, 68'b01001100101001101001101111000001100010111000110011001011010000111001); #20
	MCMC_indirect_write(11'd1142, 68'b00010101011001111001110000101001100010011001111110000011110000100010); #20
	MCMC_indirect_write(11'd1143, 68'b00111100100101011010010101100010000010101100110010000000010100010000); #20
	MCMC_indirect_write(11'd1144, 68'b01101100010110010011010000001111010110001100001010001110011000001110); #20
	MCMC_indirect_write(11'd1145, 68'b01010101101011110010001010100001000100010000101000101010111011001111); #20
	MCMC_indirect_write(11'd1146, 68'b10001111101000100101111111001100111011110010100111010110110111011100); #20
	MCMC_indirect_write(11'd1147, 68'b00010101000100110001010100111100010101001010100101000111000100001000); #20
	MCMC_indirect_write(11'd1148, 68'b11010111001100110110001011100111011011010001101001110100111011011110); #20
	MCMC_indirect_write(11'd1149, 68'b00001110111011011001011111100010100000100010100110100001000111101111); #20
	MCMC_indirect_write(11'd1150, 68'b01000011101101010010110000110101110100001101110000100110001111101000); #20
	MCMC_indirect_write(11'd1151, 68'b11010100000110101110100000111001001101101000001000010111111001101100); #20
	MCMC_indirect_write(11'd1152, 68'b10010000000000000100100000000000001001000000000000010010000000000000); #20
	MCMC_indirect_write(11'd1153, 68'b10001110101100111100100000011100010111111101100001010000001010000100); #20
	MCMC_indirect_write(11'd1154, 68'b10100110000001001100101110111011111000100000011010010001000000111100); #20
	MCMC_indirect_write(11'd1155, 68'b10111011011111110101011000100110101011110111110011010011001101100110); #20
	MCMC_indirect_write(11'd1156, 68'b10101101001010100101100000010100101010100010001000110000011011001111); #20
	MCMC_indirect_write(11'd1157, 68'b10111101000010111110101010011100101111000001101101111011000010010100); #20
	MCMC_indirect_write(11'd1158, 68'b10000000101011101100011111000111101001011110000011010100011110001011); #20
	MCMC_indirect_write(11'd1159, 68'b00110010111001111001010000100100110010100101000010101010000011111000); #20
	MCMC_indirect_write(11'd1160, 68'b01010110001001101001110101100100000100111011101011100110000000110011); #20
	MCMC_indirect_write(11'd1161, 68'b11100011111111000111011000011011110000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1162, 68'b10011011000101100101110010100101001101001101001011011001011101000111); #20
	MCMC_indirect_write(11'd1163, 68'b10100000100000101101110001010101001100000111100110010110010000000111); #20
	MCMC_indirect_write(11'd1164, 68'b11001110100001010100100110000110101010110011110101010011000101101011); #20
	MCMC_indirect_write(11'd1165, 68'b10110100000111100101111000100111101001101010110010010100110010011111); #20
	MCMC_indirect_write(11'd1166, 68'b10110001100100011101011000010100001100001100111001011010110101100010); #20
	MCMC_indirect_write(11'd1167, 68'b01011000100101101100110011100111111010010011110111010110001101000000); #20
	MCMC_indirect_write(11'd1168, 68'b00111101110110001000001000100010010000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1169, 68'b10000111111110000100111111010000111010010001111110101111100101110100); #20
	MCMC_indirect_write(11'd1170, 68'b10010100001111110011011000010001100110110100100101010011111010111110); #20
	MCMC_indirect_write(11'd1171, 68'b10110110001111111101011110111001101010011111100101111011010000111001); #20
	MCMC_indirect_write(11'd1172, 68'b10001011101111010100100101001111110111000000101010010011101000010101); #20
	MCMC_indirect_write(11'd1173, 68'b10101001010000101100100011011000001000110111110100110011010001010001); #20
	MCMC_indirect_write(11'd1174, 68'b10011101100001101110111100001111101110010000100010010000000000000000); #20
	MCMC_indirect_write(11'd1175, 68'b00110011111110010010011100000000000011100010101101000110111110010101); #20
	MCMC_indirect_write(11'd1176, 68'b10100010001110010101000101101110111100011011101101010110001101000111); #20
	MCMC_indirect_write(11'd1177, 68'b00100100000100100001011100111001100010111001011111100111101010100111); #20
	MCMC_indirect_write(11'd1178, 68'b00000110100000010000010100110000100000101100100111000010101111011000); #20
	MCMC_indirect_write(11'd1179, 68'b01101011110100000011111111111110010111001001110110010001101101110011); #20
	MCMC_indirect_write(11'd1180, 68'b11110110100100101100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1181, 68'b01111110000100010011101111011110001000100111011001001101011010000111); #20
	MCMC_indirect_write(11'd1182, 68'b01111110001111011100000001110001011000100000101011110111001111101000); #20
	MCMC_indirect_write(11'd1183, 68'b10000010010000010010111000001111010101100101001111001101011011110101); #20
	MCMC_indirect_write(11'd1184, 68'b11010110011101011110001111111111101011010010110000110111001000111100); #20
	MCMC_indirect_write(11'd1185, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1186, 68'b01011010000000101010110110110100110101100110111000001111010001010011); #20
	MCMC_indirect_write(11'd1187, 68'b01001100000001001010011010000110100110110001111101110001001011110011); #20
	MCMC_indirect_write(11'd1188, 68'b01110110100111101011010010011101110111000100001111101010100010111100); #20
	MCMC_indirect_write(11'd1189, 68'b01100001101000110011000000100111100101011001101111101110001001101101); #20
	MCMC_indirect_write(11'd1190, 68'b10010010110111100101101000100110111001011011111100010100110000100101); #20
	MCMC_indirect_write(11'd1191, 68'b10100011011101100101010000101110001001010001011100110011110111100101); #20
	MCMC_indirect_write(11'd1192, 68'b11010100001010100100000000000000001111100100101100111001110000000101); #20
	MCMC_indirect_write(11'd1193, 68'b10111111111100100110010001000100101011111011001111111011100010100001); #20
	MCMC_indirect_write(11'd1194, 68'b10010010001111101011100001110000100101001001110010001011000011111011); #20
	MCMC_indirect_write(11'd1195, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1196, 68'b11101110011011011100000000000000001000000000000000011110101111011110); #20
	MCMC_indirect_write(11'd1197, 68'b01111100100010100010010101100001110110010110101000101011000001110011); #20
	MCMC_indirect_write(11'd1198, 68'b11100110000101100111001011110101001101011001111000110111010100011011); #20
	MCMC_indirect_write(11'd1199, 68'b10101001000010110101111100000010111011101000111111111101000110010101); #20
	MCMC_indirect_write(11'd1200, 68'b10000000000000000011110101010011000111000101001001111011110010000111); #20
	MCMC_indirect_write(11'd1201, 68'b10101100000111011101101010101000111010100011101111010110000001100100); #20
	MCMC_indirect_write(11'd1202, 68'b11000100111100101110110000000000001110000001000110010000000000000000); #20
	MCMC_indirect_write(11'd1203, 68'b11000101011011000101110011000111011000110000111010110000000100111110); #20
	MCMC_indirect_write(11'd1204, 68'b00011100100010111001011001101010010100000110111111100101101010011111); #20
	MCMC_indirect_write(11'd1205, 68'b01010101011000111010010111001110110100011000101000101000001010010111); #20
	MCMC_indirect_write(11'd1206, 68'b10101010010010011100111110001011111011000000011110110101010101011011); #20
	MCMC_indirect_write(11'd1207, 68'b10010100011111000101010000001011001011100001101110011010110000001110); #20
	MCMC_indirect_write(11'd1208, 68'b11010011010000110110100000000100011101110110110011011011110001100000); #20
	MCMC_indirect_write(11'd1209, 68'b10001010010001010010010000000100100101111001010100001110111111011110); #20
	MCMC_indirect_write(11'd1210, 68'b01010110000100001011000101000101000011111111011110100000110110011110); #20
	MCMC_indirect_write(11'd1211, 68'b11011111111011110110011011100000001011111110001010110101000000010010); #20
	MCMC_indirect_write(11'd1212, 68'b11011010100101001111100011000000001101010110101000011011111101101111); #20
	MCMC_indirect_write(11'd1213, 68'b10010000101000010101111111101011111110101011101010110000000000000000); #20
	MCMC_indirect_write(11'd1214, 68'b01010010100100001001010110011010000011111111110010000110000001001100); #20
	MCMC_indirect_write(11'd1215, 68'b10111101010110010101110000001010111011000101010001110011110001110001); #20
	MCMC_indirect_write(11'd1216, 68'b10011000000000000100110000000000001001100000000000010011000000000000); #20
	MCMC_indirect_write(11'd1217, 68'b10001100001111010100000001110110101000011000111010010100100101110001); #20
	MCMC_indirect_write(11'd1218, 68'b10010000111001011100110110010000111011000010100011010010110100111011); #20
	MCMC_indirect_write(11'd1219, 68'b10100110100111011100000000010110111000100100010000010010101111000001); #20
	MCMC_indirect_write(11'd1220, 68'b10100110110111100100010010100101111010000001100100001111101100111000); #20
	MCMC_indirect_write(11'd1221, 68'b01100011010101101010111001100001110101111011010010001101000101110001); #20
	MCMC_indirect_write(11'd1222, 68'b11001110000110001100111011110111000111001100011110101011111001000101); #20
	MCMC_indirect_write(11'd1223, 68'b11010100100001101110110010001100101011110001001101111010110011000111); #20
	MCMC_indirect_write(11'd1224, 68'b10011010110011000100111010101101001000101111011101110010100101001100); #20
	MCMC_indirect_write(11'd1225, 68'b11010000110011110101101111011111001011101111111000011111000110100000); #20
	MCMC_indirect_write(11'd1226, 68'b01110011100010111100000111000011001000110101101110110000000101001011); #20
	MCMC_indirect_write(11'd1227, 68'b01001110001111101010101001010010100110111111100001100101101001110001); #20
	MCMC_indirect_write(11'd1228, 68'b11101100000010111101011010101111101010010000110100110011010001001001); #20
	MCMC_indirect_write(11'd1229, 68'b00100110110101101010011001100000000100111000100011001000000111101110); #20
	MCMC_indirect_write(11'd1230, 68'b10100110101010000100100000110110111100001010101001010110011001001111); #20
	MCMC_indirect_write(11'd1231, 68'b10111100110011101110010111100100111100011011111100111011001001001000); #20
	MCMC_indirect_write(11'd1232, 68'b10000011001100010011111001010110000110011100101011010000100011100110); #20
	MCMC_indirect_write(11'd1233, 68'b01110100100101011011101011001100011000111011000110010100000001000100); #20
	MCMC_indirect_write(11'd1234, 68'b10000000110101110100100100110010001010100011110000010000011001001011); #20
	MCMC_indirect_write(11'd1235, 68'b10001000000111101101011001000100111011100101110000110010010111000101); #20
	MCMC_indirect_write(11'd1236, 68'b00111010110111110010100110111100010100100101010010100110100000010000); #20
	MCMC_indirect_write(11'd1237, 68'b10101000110111011101100001000100011011100101011111110100010101101110); #20
	MCMC_indirect_write(11'd1238, 68'b10011111010100111110000100001011101011101001010011110110100110111101); #20
	MCMC_indirect_write(11'd1239, 68'b11110111011100101111001111001011101101000000001000010111100000110001); #20
	MCMC_indirect_write(11'd1240, 68'b01100100110011100011001110011000000101110100000011101100111000100110); #20
	MCMC_indirect_write(11'd1241, 68'b10000000000000000100000000000000010000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1242, 68'b01000000110101110001111101110111010100011000000001100111010111110011); #20
	MCMC_indirect_write(11'd1243, 68'b10010010100001010100011001100011100101100000101100001010000100010010); #20
	MCMC_indirect_write(11'd1244, 68'b01000011110100011000101000010101000001000001000001100001010101100101); #20
	MCMC_indirect_write(11'd1245, 68'b01110011110111011011110110101011011001000100111101010100100001110111); #20
	MCMC_indirect_write(11'd1246, 68'b01101100110001110100010011100010111011100010011000010110011101110001); #20
	MCMC_indirect_write(11'd1247, 68'b01101000000000110011100000110010011001000010110001010000100101100000); #20
	MCMC_indirect_write(11'd1248, 68'b00111000100111000001111001101010000010001000001110100010101010001011); #20
	MCMC_indirect_write(11'd1249, 68'b10000011010011110101100101111110011011111111111110011000001101110101); #20
	MCMC_indirect_write(11'd1250, 68'b11000101000101110110011001011000011110001101110001010111110000010000); #20
	MCMC_indirect_write(11'd1251, 68'b01111100001010010010110110111101110100111010110000101011111110000110); #20
	MCMC_indirect_write(11'd1252, 68'b00111110010100011010010011110101110110110101001100110001001110011111); #20
	MCMC_indirect_write(11'd1253, 68'b01110000101001001100001110001110111000100100101011001110111011010100); #20
	MCMC_indirect_write(11'd1254, 68'b01000110110001110011001111101011110100000000010111000110110011011100); #20
	MCMC_indirect_write(11'd1255, 68'b01010011001101111001001100110111010001110101000100000011111000001100); #20
	MCMC_indirect_write(11'd1256, 68'b10000101100001011011100000000110110110011011010100000110010001010100); #20
	MCMC_indirect_write(11'd1257, 68'b11010110101011010110001010110110001001010000000101011000001001001010); #20
	MCMC_indirect_write(11'd1258, 68'b00010111100111001000111100111011100001001101011001101000101111101101); #20
	MCMC_indirect_write(11'd1259, 68'b10010100010011101101101001111110111110000010011110111011111000000101); #20
	MCMC_indirect_write(11'd1260, 68'b01010000000111011010100010110000100011001101100111001000000000000110); #20
	MCMC_indirect_write(11'd1261, 68'b10111100011010100100111001010010001010010001111100110111011000000101); #20
	MCMC_indirect_write(11'd1262, 68'b00110000101001010001010000000100000000111011110010000000010010111100); #20
	MCMC_indirect_write(11'd1263, 68'b01111001010101000011001110111001110111111101001111010001010110001001); #20
	MCMC_indirect_write(11'd1264, 68'b00000000000000000001011101001000000011110010101001100111111100001110); #20
	MCMC_indirect_write(11'd1265, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1266, 68'b11100001010111111110111001001011001111010010111101010000000000000000); #20
	MCMC_indirect_write(11'd1267, 68'b01000101000000000001001101010110100000000001010001000001010101010011); #20
	MCMC_indirect_write(11'd1268, 68'b10110110001100101101100110110100011001111101001000110011001101101101); #20
	MCMC_indirect_write(11'd1269, 68'b01111100000011001100011000111010101001011110000101010010010110001000); #20
	MCMC_indirect_write(11'd1270, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1271, 68'b10111100100111010101100000011110101000011101000011010001000101101001); #20
	MCMC_indirect_write(11'd1272, 68'b00000010010100010000000000000000000001011100001000000110011001111110); #20
	MCMC_indirect_write(11'd1273, 68'b11010001101001101101101111011100111010001011100110010100111111000011); #20
	MCMC_indirect_write(11'd1274, 68'b10011000011100000011010001011101100111001101010001010000110001001000); #20
	MCMC_indirect_write(11'd1275, 68'b01101110010100111011111011010100110111101011000100101101010000000110); #20
	MCMC_indirect_write(11'd1276, 68'b11101100011011111110111100001111001111000100000000100000000000000000); #20
	MCMC_indirect_write(11'd1277, 68'b10111001111110010101010111110101111001101011101010110000000100111110); #20
	MCMC_indirect_write(11'd1278, 68'b00101110100001110010100010011010000011010011110010000010011010011101); #20
	MCMC_indirect_write(11'd1279, 68'b11101101100000011111110011010111111000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1280, 68'b10100000000000000101000000000000001010000000000000010100000000000000); #20
	MCMC_indirect_write(11'd1281, 68'b10010111111001110101000000001011011001011111011111010011010000000010); #20
	MCMC_indirect_write(11'd1282, 68'b10100011100101011100001111000110101001101000111110110110010001011011); #20
	MCMC_indirect_write(11'd1283, 68'b10000001001011011100110010001100001001010110001100110000000001010101); #20
	MCMC_indirect_write(11'd1284, 68'b10100110010001001100111100110010101011110100000111010110100100000101); #20
	MCMC_indirect_write(11'd1285, 68'b10111110000111011100101010101111111001101000011111010110111000101011); #20
	MCMC_indirect_write(11'd1286, 68'b00110100001100010001011011010101100010111011000110001000100100011010); #20
	MCMC_indirect_write(11'd1287, 68'b10001011101011010100001100001011111010101001110000010011000110001010); #20
	MCMC_indirect_write(11'd1288, 68'b10001110000000000101100101011100001001110110010110111001101101111001); #20
	MCMC_indirect_write(11'd1289, 68'b10000000000000000100000000000000001101001101111110111001101101001110); #20
	MCMC_indirect_write(11'd1290, 68'b01001100111001001010010010000110100100110000000100101010101111100000); #20
	MCMC_indirect_write(11'd1291, 68'b01010011001001001010110010110010110100010100011010101001001110110001); #20
	MCMC_indirect_write(11'd1292, 68'b01110011010101001010111101011001000011011011001000100011000100101011); #20
	MCMC_indirect_write(11'd1293, 68'b10111011001010011101010000011001011011010010010101010110011011101101); #20
	MCMC_indirect_write(11'd1294, 68'b10000110011101000110000001010001111011101011111110010111101001011101); #20
	MCMC_indirect_write(11'd1295, 68'b11010100011100000111011011101001111110110011100001011000100101000100); #20
	MCMC_indirect_write(11'd1296, 68'b10001100010000110100001000111100001000100000110110001101111010011101); #20
	MCMC_indirect_write(11'd1297, 68'b01101000110011111010111111100000000111110110101011101110011000111001); #20
	MCMC_indirect_write(11'd1298, 68'b10101000110111100110001111100000011101101011011100111011011010000111); #20
	MCMC_indirect_write(11'd1299, 68'b10011110101000001100110000111011101000110010111101110110010110011110); #20
	MCMC_indirect_write(11'd1300, 68'b10101100001010100100110111011011001011100001100000010000111110000011); #20
	MCMC_indirect_write(11'd1301, 68'b01010111001001100011111110111001110111101111000110110010010110111111); #20
	MCMC_indirect_write(11'd1302, 68'b11011000111101001110001100001010011001110001110001110101001000011010); #20
	MCMC_indirect_write(11'd1303, 68'b01100111011011001100010111000100110111101010110011110001001100110101); #20
	MCMC_indirect_write(11'd1304, 68'b11101011111001011111010001110011011100010011011111100000000000000000); #20
	MCMC_indirect_write(11'd1305, 68'b11011000010000010111000000001011011011101111000000110001111110101000); #20
	MCMC_indirect_write(11'd1306, 68'b10010001011010111100011011001011011001100011101010110011010011010010); #20
	MCMC_indirect_write(11'd1307, 68'b10001001001110110010111100001000010111000011111011001110100101011101); #20
	MCMC_indirect_write(11'd1308, 68'b00000000000101111000110001001001110001100001111010100000000000000000); #20
	MCMC_indirect_write(11'd1309, 68'b10011110011010110100010001001001110101000110101011000011111000110111); #20
	MCMC_indirect_write(11'd1310, 68'b11000011111001111110101111010001110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1311, 68'b10000000000000000111100100111010110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1312, 68'b01101100111010001001111101111011100011011001100010000110010010011010); #20
	MCMC_indirect_write(11'd1313, 68'b10100011111101100101101100101011111011111011111100110111110111110000); #20
	MCMC_indirect_write(11'd1314, 68'b01011001010011010010011000101101010100110000000110001100000110011010); #20
	MCMC_indirect_write(11'd1315, 68'b10100001011111010100111111110110111000011010011010010001100100000101); #20
	MCMC_indirect_write(11'd1316, 68'b10000111110100100100001001011001110111101100111010110010110011001010); #20
	MCMC_indirect_write(11'd1317, 68'b11100111101110001111010110101100001110101111011011111110010110101001); #20
	MCMC_indirect_write(11'd1318, 68'b10110101101110110101110100110111001011110000011011011100011101011100); #20
	MCMC_indirect_write(11'd1319, 68'b01111010101111101011011000000010010111101010100100001111110101100001); #20
	MCMC_indirect_write(11'd1320, 68'b01111110110011001011100101000110110111111010011101010101011001011100); #20
	MCMC_indirect_write(11'd1321, 68'b00110101011000001010101111101101000101100011001101101100101110111001); #20
	MCMC_indirect_write(11'd1322, 68'b10000000000000000011110111100001011110001100100111111100100101111100); #20
	MCMC_indirect_write(11'd1323, 68'b10000001110101110100101110111111101011000111010000011000100100111010); #20
	MCMC_indirect_write(11'd1324, 68'b10000000000000001111011001100111010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1325, 68'b00100011001001010001010011011110010001101111110111000100011010101011); #20
	MCMC_indirect_write(11'd1326, 68'b10101101101010110110101001011000101110110100000110110000000000000000); #20
	MCMC_indirect_write(11'd1327, 68'b00011111011010001000101000111000010000000000000000000000110101111011); #20
	MCMC_indirect_write(11'd1328, 68'b01011101110110101010101000110000110110011011010010010000100111110000); #20
	MCMC_indirect_write(11'd1329, 68'b00110010101010010001101000110010010100011000110101100011100010000111); #20
	MCMC_indirect_write(11'd1330, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1331, 68'b10010101000001110110101001110011111101101011000101011000101000101011); #20
	MCMC_indirect_write(11'd1332, 68'b10000101111100101100100111101110001001111100000100110011101001001001); #20
	MCMC_indirect_write(11'd1333, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1334, 68'b11100011001011010101111111010001101010010100000011010110011011000011); #20
	MCMC_indirect_write(11'd1335, 68'b10101111011010111100110011001110011010011011001100111001110101111100); #20
	MCMC_indirect_write(11'd1336, 68'b01011010000111110011010111110101111011010101111100010001011001010001); #20
	MCMC_indirect_write(11'd1337, 68'b11110111100101001111011001001101001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1338, 68'b10101000011101111100001111010110111001101100101011110011000101100011); #20
	MCMC_indirect_write(11'd1339, 68'b10000000000000000010000000000000000100000000000000001110011011010101); #20
	MCMC_indirect_write(11'd1340, 68'b11010111101001011111101010110110010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1341, 68'b01010110010011110010101000010110110011001110110000100110010010011100); #20
	MCMC_indirect_write(11'd1342, 68'b10010100110010011011011111001010011001001010110011001011011011011111); #20
	MCMC_indirect_write(11'd1343, 68'b10100100101001101100011010001011111010110110101001010010100000110011); #20
	MCMC_indirect_write(11'd1344, 68'b10101000000000000101010000000000001010100000000000010101000000000000); #20
	MCMC_indirect_write(11'd1345, 68'b10101000110101011101011000111010101010100001101011110100111100110011); #20
	MCMC_indirect_write(11'd1346, 68'b10100100011000010101111110111111101000111111010010110010000001011101); #20
	MCMC_indirect_write(11'd1347, 68'b10001000010100011100011111000100101010001010010010010001111001011010); #20
	MCMC_indirect_write(11'd1348, 68'b10010100100110001101001100100010101001011011001111110111101000101100); #20
	MCMC_indirect_write(11'd1349, 68'b01110010001011101001111000010000010011110001010100101000111010011110); #20
	MCMC_indirect_write(11'd1350, 68'b10001111011110111100000101101100110100010111000101101100100001100111); #20
	MCMC_indirect_write(11'd1351, 68'b11011000110011001111001000111000110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1352, 68'b01101111110010110100000100010001011000011100010010010001000001010000); #20
	MCMC_indirect_write(11'd1353, 68'b10100011110011001101010110101000111100111011111011110011010010111101); #20
	MCMC_indirect_write(11'd1354, 68'b11101001001010111100000000000000001000000000000000011101101111011101); #20
	MCMC_indirect_write(11'd1355, 68'b11101110000101001110001001101101110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1356, 68'b00110100110111001001100011111011010001110010010001100001110110110001); #20
	MCMC_indirect_write(11'd1357, 68'b10000010010010111100001100100110001000101000110110110010000001010001); #20
	MCMC_indirect_write(11'd1358, 68'b11000010110011000110010011110011011100011011011110110000000000000000); #20
	MCMC_indirect_write(11'd1359, 68'b10000000000000000010000000000000000100000000000000001000000000000000); #20
	MCMC_indirect_write(11'd1360, 68'b11011111000111000110101010000000011100101100010111010100110000111011); #20
	MCMC_indirect_write(11'd1361, 68'b11011101111110010110110011110010111101000001010101010101111011101001); #20
	MCMC_indirect_write(11'd1362, 68'b11001110011010001101111110110000001110001100101110011111001010100011); #20
	MCMC_indirect_write(11'd1363, 68'b11010001010011110101110000001110101011011111010100010111111111010100); #20
	MCMC_indirect_write(11'd1364, 68'b11000011000001100110011100100100111101110111001011110111010111101010); #20
	MCMC_indirect_write(11'd1365, 68'b00110001111100111001000111000000000001011011011101101000001101100111); #20
	MCMC_indirect_write(11'd1366, 68'b10100000000100101011100101000100000101111011000011100110011111010110); #20
	MCMC_indirect_write(11'd1367, 68'b10100001111111010100100001000100011001110111001010010111110011111111); #20
	MCMC_indirect_write(11'd1368, 68'b01100000010110011011000011011011100011111110111000000111100010011000); #20
	MCMC_indirect_write(11'd1369, 68'b10010110100111001100000011011100001000011001001101010000111100000000); #20
	MCMC_indirect_write(11'd1370, 68'b10000000000000000011111000000011010111100011110101011010111110011111); #20
	MCMC_indirect_write(11'd1371, 68'b11001111001010111101101010010110111101010101110000100000000000000000); #20
	MCMC_indirect_write(11'd1372, 68'b01010100110000110011011001000101110101000010111001101110011000010110); #20
	MCMC_indirect_write(11'd1373, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1374, 68'b10100001011101100101100011100011101000100100011100110001000001111000); #20
	MCMC_indirect_write(11'd1375, 68'b00110111010110000010100000010101100000111100100100000000000000000000); #20
	MCMC_indirect_write(11'd1376, 68'b11110100101101111111000100010011101100010000100011001111101101000001); #20
	MCMC_indirect_write(11'd1377, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1378, 68'b01011001101010110011010111000100100101011000110101101000110110100111); #20
	MCMC_indirect_write(11'd1379, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1380, 68'b10101110000010001011111111111010101000111011011001110110111100110010); #20
	MCMC_indirect_write(11'd1381, 68'b01101100110100000010100010000011000101001010101111101001110010101011); #20
	MCMC_indirect_write(11'd1382, 68'b01101001110110011010110000001001010011111000000010000101000010001111); #20
	MCMC_indirect_write(11'd1383, 68'b11000010110011101110101101010001111110010010100011111000011011100000); #20
	MCMC_indirect_write(11'd1384, 68'b01111001110101010010011111000100100111100011000001101111011011001011); #20
	MCMC_indirect_write(11'd1385, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1386, 68'b00110100101110111001100010111011110011011101101110101100100000101100); #20
	MCMC_indirect_write(11'd1387, 68'b10011111000001001100110001100100111010011100000100110100011111000011); #20
	MCMC_indirect_write(11'd1388, 68'b10011101101100000110001100111010011010111110000100110111010011000000); #20
	MCMC_indirect_write(11'd1389, 68'b01011111111010100010101000110111100100110011001101101010000010110011); #20
	MCMC_indirect_write(11'd1390, 68'b11100101010110111011111011100111011010100111101110100000000000000000); #20
	MCMC_indirect_write(11'd1391, 68'b10000000000000000100000000000000001000000000000000011101101001100010); #20
	MCMC_indirect_write(11'd1392, 68'b10110101100001000101001001011110011011001001110110111000011111011000); #20
	MCMC_indirect_write(11'd1393, 68'b10010000011100101100000111001110010110001101011100010001011011010111); #20
	MCMC_indirect_write(11'd1394, 68'b00011110000000110000101110011110010001101000001101000101011010100001); #20
	MCMC_indirect_write(11'd1395, 68'b01111011110110011011010000001111010110111010001010010011100011111001); #20
	MCMC_indirect_write(11'd1396, 68'b10011001111100010011110010000001000111011011110101110100000110011110); #20
	MCMC_indirect_write(11'd1397, 68'b10000000000000000111001000100010011100010010010001010111100001110111); #20
	MCMC_indirect_write(11'd1398, 68'b11100011101100111111010101000000011101100001100110010111011101001101); #20
	MCMC_indirect_write(11'd1399, 68'b11101111111011110110010101010111001100011111001110110101000011000000); #20
	MCMC_indirect_write(11'd1400, 68'b01001011111010111010110100001101110100010111101011000111011111110010); #20
	MCMC_indirect_write(11'd1401, 68'b11000101110111001101111000001010001010000001011101110110100000000001); #20
	MCMC_indirect_write(11'd1402, 68'b10001101100110000100011110010001111001011100001011110001100011011000); #20
	MCMC_indirect_write(11'd1403, 68'b10100010010000111100100010001010011001001101110100001111000011011011); #20
	MCMC_indirect_write(11'd1404, 68'b01100100000100100010010001100001110101101101110000101100100100111011); #20
	MCMC_indirect_write(11'd1405, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1406, 68'b00101111000101101010101001100011100101010001100010001110010010010000); #20
	MCMC_indirect_write(11'd1407, 68'b10011110110111010101000001100110001011111100111001010111001111100011); #20
	MCMC_indirect_write(11'd1408, 68'b10110000000000000101100000000000001011000000000000010110000000000000); #20
	MCMC_indirect_write(11'd1409, 68'b10110001101100101101010101001001101010100100111110110110100010010110); #20
	MCMC_indirect_write(11'd1410, 68'b10001111010100100110011000110111011100011100010010010100010110010110); #20
	MCMC_indirect_write(11'd1411, 68'b10101100010010100101001010111000101010100100101101010110101100010101); #20
	MCMC_indirect_write(11'd1412, 68'b10101101101011100100110110011001011010001111010111110101011100100010); #20
	MCMC_indirect_write(11'd1413, 68'b10101101111101010110101000110001001100101010010010110111100101101011); #20
	MCMC_indirect_write(11'd1414, 68'b10000111001111101011101111001000010110100000100111001101110111000000); #20
	MCMC_indirect_write(11'd1415, 68'b10100101011000101110000010110101111011010111011110010110100100010001); #20
	MCMC_indirect_write(11'd1416, 68'b10101110111101111100110011000010001001110001110100011001101000010101); #20
	MCMC_indirect_write(11'd1417, 68'b10110101001010001101111000100100111100110100001111011100101111100110); #20
	MCMC_indirect_write(11'd1418, 68'b01110110010100111100010100001100111011011001110101011001001000001111); #20
	MCMC_indirect_write(11'd1419, 68'b10011100011110010011111001010010111000000110010001010000010011100011); #20
	MCMC_indirect_write(11'd1420, 68'b01110101100101000011101110100011110110001110100111001101011100101010); #20
	MCMC_indirect_write(11'd1421, 68'b00011110010000111001010000011010010011001000101100100110100000100010); #20
	MCMC_indirect_write(11'd1422, 68'b10110011100111111110111000010000101110010000100101011110111000010111); #20
	MCMC_indirect_write(11'd1423, 68'b01000001100011110000111101000001000100000100100000001100001111101010); #20
	MCMC_indirect_write(11'd1424, 68'b10111000111110001101000100101001001001111101001011010110011110100000); #20
	MCMC_indirect_write(11'd1425, 68'b00110000011110011001010010001010110100001010111011000011011010011100); #20
	MCMC_indirect_write(11'd1426, 68'b10000000000000000011111011011110010111000010000011101010011011010101); #20
	MCMC_indirect_write(11'd1427, 68'b01110000100110010100000011100111100110100100101101001100001000101100); #20
	MCMC_indirect_write(11'd1428, 68'b10001011011011010100111101001101111001001110110011001100111100100001); #20
	MCMC_indirect_write(11'd1429, 68'b00111010110110010001101111100010110001100110000100100100011101111101); #20
	MCMC_indirect_write(11'd1430, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1431, 68'b10001101000010101100111101111111011001111000001010110110001011011011); #20
	MCMC_indirect_write(11'd1432, 68'b11000101010111000101001111110100011100000000101101010111011001000111); #20
	MCMC_indirect_write(11'd1433, 68'b01110101110010010011111011010110110110111010100000001110000100000011); #20
	MCMC_indirect_write(11'd1434, 68'b11110011111110111110001101101000110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1435, 68'b10000000000000000010000000000000000111001111100101111011111000110000); #20
	MCMC_indirect_write(11'd1436, 68'b01110101000001101010011110000001010100101100111001000101000111100010); #20
	MCMC_indirect_write(11'd1437, 68'b01011001101111100010100101111111100011110101111110101000101110101001); #20
	MCMC_indirect_write(11'd1438, 68'b00111011101000011011011000100001010101001000110111001011101001010111); #20
	MCMC_indirect_write(11'd1439, 68'b01110100011000100101010100010111001100100000011010110110011100110110); #20
	MCMC_indirect_write(11'd1440, 68'b10001110100001100011111000101101100110100110100000001001101000011110); #20
	MCMC_indirect_write(11'd1441, 68'b11000001001111110111010101110101011000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1442, 68'b01111101000110101011111101011101010111001110100111110001011101011010); #20
	MCMC_indirect_write(11'd1443, 68'b10000000101110111011001110110111000101111100011100110000000010100001); #20
	MCMC_indirect_write(11'd1444, 68'b11111000010111011100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1445, 68'b10111111000010111110001010001011001011101011010111110111100010111010); #20
	MCMC_indirect_write(11'd1446, 68'b10010000010001010100000110101111010111010001110101101100011011100100); #20
	MCMC_indirect_write(11'd1447, 68'b10100001101000000100010110111110011001111101010010010110010101100110); #20
	MCMC_indirect_write(11'd1448, 68'b10010111110001000101111111101111001100100100101011110011111000011111); #20
	MCMC_indirect_write(11'd1449, 68'b11011111011110100101010111000111011010100000010010010110110100101110); #20
	MCMC_indirect_write(11'd1450, 68'b11101100110100101111101011011101011000000000000000011101001100100011); #20
	MCMC_indirect_write(11'd1451, 68'b10011111010001111100111011111011001001001101111001010011110010111000); #20
	MCMC_indirect_write(11'd1452, 68'b11101110011111111111110011010100011111110111100000011110101010101110); #20
	MCMC_indirect_write(11'd1453, 68'b10101111110101110101000100000010111001001110110100011010010001000001); #20
	MCMC_indirect_write(11'd1454, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1455, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1456, 68'b11011011101001010111010011011100111101010111100001011010110110001111); #20
	MCMC_indirect_write(11'd1457, 68'b10101000000100001100001001001110010101111101110010101100111001110000); #20
	MCMC_indirect_write(11'd1458, 68'b10100011111010111100110000101111101011100110000101111001110101110100); #20
	MCMC_indirect_write(11'd1459, 68'b11110011111110011111110100000110010000000000000000011100010011111001); #20
	MCMC_indirect_write(11'd1460, 68'b11101101000101100110111010001000011100110010100001011100111000010001); #20
	MCMC_indirect_write(11'd1461, 68'b11100100011111001111110110100101110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1462, 68'b01001000001010100001100110010101110010111100110011100101110011010110); #20
	MCMC_indirect_write(11'd1463, 68'b01100100000110110010100010001000110100011011000111000111101111011001); #20
	MCMC_indirect_write(11'd1464, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1465, 68'b11000011010010100110011001000100011011001001100000110101100000000000); #20
	MCMC_indirect_write(11'd1466, 68'b10010000100011001100010001011100011000101011011010010000011100001111); #20
	MCMC_indirect_write(11'd1467, 68'b11011101011111011111001011011110010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1468, 68'b00111011110010110001100110011100100010100011111000100111000011001101); #20
	MCMC_indirect_write(11'd1469, 68'b11001101100101101110001111000010111101000011110111011011010011101011); #20
	MCMC_indirect_write(11'd1470, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1471, 68'b11010101110001111110001010010110001011101001110111010110111111110100); #20
	MCMC_indirect_write(11'd1472, 68'b10111000000000000101110000000000001011100000000000010111000000000000); #20
	MCMC_indirect_write(11'd1473, 68'b10110011100001011101111001110001001011010100011001110110111000000000); #20
	MCMC_indirect_write(11'd1474, 68'b10101001011100000110001001101101011010001000100011110110100101010000); #20
	MCMC_indirect_write(11'd1475, 68'b10110110000010000110001010110001001100101100011101011100011111011100); #20
	MCMC_indirect_write(11'd1476, 68'b11000000110110101110000101011011101010110100110011110111011111011110); #20
	MCMC_indirect_write(11'd1477, 68'b10000001110010000100100100111100101011101111001010111000010111001111); #20
	MCMC_indirect_write(11'd1478, 68'b10110111000110111110100011001000001100011010100001111100111010101000); #20
	MCMC_indirect_write(11'd1479, 68'b11010100100001100101101010101100101011101100110110110110001010110101); #20
	MCMC_indirect_write(11'd1480, 68'b11010101101010111110111011000011001100001001000100011000010100010111); #20
	MCMC_indirect_write(11'd1481, 68'b11111010100011000111110011100001001100001101101000111000000011101000); #20
	MCMC_indirect_write(11'd1482, 68'b11111010101000000100000000000000001000000000000000011101010101011100); #20
	MCMC_indirect_write(11'd1483, 68'b10110101110000011101101101110111111010010101101100010010001010100000); #20
	MCMC_indirect_write(11'd1484, 68'b11000111110111101101110001101010111001111001101101010011111011101011); #20
	MCMC_indirect_write(11'd1485, 68'b01111001000000010011110010111100000110110101111110001100110001011111); #20
	MCMC_indirect_write(11'd1486, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1487, 68'b10000110000110110110000101111010011001011011001101010101011011011100); #20
	MCMC_indirect_write(11'd1488, 68'b11001100011110000110101000010011101110101100101011111101100111100111); #20
	MCMC_indirect_write(11'd1489, 68'b10000000000000000111010100010011001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1490, 68'b10110110000001001110011101011111101010111110001001011001111110001011); #20
	MCMC_indirect_write(11'd1491, 68'b11100110001101111111011010000010101111000110110101011101011001101110); #20
	MCMC_indirect_write(11'd1492, 68'b11011001000100100111000111101110001101001011011111110111111011111000); #20
	MCMC_indirect_write(11'd1493, 68'b10111111100101100110000111010010001000111111001101110010010100000010); #20
	MCMC_indirect_write(11'd1494, 68'b01010101100100100011011010110010111000011010001001001010100110101000); #20
	MCMC_indirect_write(11'd1495, 68'b10100110101101111101101001010001011101000110000100111000010110101100); #20
	MCMC_indirect_write(11'd1496, 68'b11000101000011000101100101011110101011011000011011110101000101000010); #20
	MCMC_indirect_write(11'd1497, 68'b10001100000001001100010110000000001001100110011000010110011101110000); #20
	MCMC_indirect_write(11'd1498, 68'b01101100111010010010110011101111000011100001111011101100111100100010); #20
	MCMC_indirect_write(11'd1499, 68'b10000000000000000011111001100010111110111101000101101100111010000010); #20
	MCMC_indirect_write(11'd1500, 68'b01010001110010100001100101110000010001110010000000100010011100101010); #20
	MCMC_indirect_write(11'd1501, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1502, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1503, 68'b11000110110001011110110001101011101110101111000110111100001000101101); #20
	MCMC_indirect_write(11'd1504, 68'b01011011111011110001111000011000010100100111100111101001011111101001); #20
	MCMC_indirect_write(11'd1505, 68'b11000001000111010101001111011100011100000010011100111000111010101001); #20
	MCMC_indirect_write(11'd1506, 68'b10011011110100110101001000100011001100000010100000111001000000101011); #20
	MCMC_indirect_write(11'd1507, 68'b10000111101011100100000101011110000111111001000101101110111001101101); #20
	MCMC_indirect_write(11'd1508, 68'b11101000011000100111010110001001010000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1509, 68'b10011100001100010101011000010010111001100100011001010000000011100011); #20
	MCMC_indirect_write(11'd1510, 68'b01111011011100110011111100010010010110010111010101001010100100100001); #20
	MCMC_indirect_write(11'd1511, 68'b01011111001111100100111100011001111001100110011000010001001001111101); #20
	MCMC_indirect_write(11'd1512, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1513, 68'b11001110100101101111101000011001111110100000100101111111100000010011); #20
	MCMC_indirect_write(11'd1514, 68'b00001000000001110001100001101011100011000010000100000010000101100110); #20
	MCMC_indirect_write(11'd1515, 68'b11001001011101001101110011001001101001100010001111110100111011001000); #20
	MCMC_indirect_write(11'd1516, 68'b10101000001110000101000011000000001010000111100100110111100010011011); #20
	MCMC_indirect_write(11'd1517, 68'b01101111111100001011000101111011100101000011010000000101011111010010); #20
	MCMC_indirect_write(11'd1518, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1519, 68'b10110100100010100011111111000110001010000011101011010010000101010111); #20
	MCMC_indirect_write(11'd1520, 68'b10100010110110101100011100010110000111101000110010010100011101011001); #20
	MCMC_indirect_write(11'd1521, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1522, 68'b11111100100100110110011111111001101011001101101011010101001111000001); #20
	MCMC_indirect_write(11'd1523, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1524, 68'b00111111111001001001110011110111110010111001010101000100010011010010); #20
	MCMC_indirect_write(11'd1525, 68'b01111110110100001011111000010010101001001100110000010010011000101011); #20
	MCMC_indirect_write(11'd1526, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1527, 68'b11001111010000001110000110010000111100001101110001110110111111100011); #20
	MCMC_indirect_write(11'd1528, 68'b11100111100011011000000000000000010000000000000000011110010011011110); #20
	MCMC_indirect_write(11'd1529, 68'b10101011110101000101001001011110011001111010111111010011001001001011); #20
	MCMC_indirect_write(11'd1530, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1531, 68'b11010110001000010110000000010001101010010110110000010011110111000010); #20
	MCMC_indirect_write(11'd1532, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1533, 68'b01011011111100101010101111111100000110001001000001001010100111010010); #20
	MCMC_indirect_write(11'd1534, 68'b01010111010110101010011111110000000001010111100111100011100111100010); #20
	MCMC_indirect_write(11'd1535, 68'b11010111111011000110001001101110101100111110101000010000000000000000); #20
	MCMC_indirect_write(11'd1536, 68'b11000000000000000110000000000000001100000000000000011000000000000000); #20
	MCMC_indirect_write(11'd1537, 68'b11000101100101001110010000100100101011011001000010011001100111110101); #20
	MCMC_indirect_write(11'd1538, 68'b11001101101111110101101001110101101100011011111011110111010010000111); #20
	MCMC_indirect_write(11'd1539, 68'b10101111010010011101101010110011111100001001111111111001110010010110); #20
	MCMC_indirect_write(11'd1540, 68'b10011000100111100100100001010010101010011001101110010111111010111001); #20
	MCMC_indirect_write(11'd1541, 68'b11001111111011011101000111110001001000110100111000010011001000010001); #20
	MCMC_indirect_write(11'd1542, 68'b01001000111000111011100010000110111000010110110110001110001001000001); #20
	MCMC_indirect_write(11'd1543, 68'b11000101010011100101101000000000101011000111101000010011100000101100); #20
	MCMC_indirect_write(11'd1544, 68'b11010101111101001101011000011010111010101110010100110110111101111110); #20
	MCMC_indirect_write(11'd1545, 68'b10110001011000001101100111100100001011101100111000111011011001100111); #20
	MCMC_indirect_write(11'd1546, 68'b01100001111110100011010100101101100110001000000010101010000101010001); #20
	MCMC_indirect_write(11'd1547, 68'b10110101110110000101101101101001101100011011000111011110101001010100); #20
	MCMC_indirect_write(11'd1548, 68'b11100010110001111111010111001100001100001000110001011001011000001000); #20
	MCMC_indirect_write(11'd1549, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1550, 68'b10100001010001100101010001101101101011001101111101010001110100000001); #20
	MCMC_indirect_write(11'd1551, 68'b00111001010010011001001010000001000010001111000100000000000000000000); #20
	MCMC_indirect_write(11'd1552, 68'b10011011010001101011110100111011111000011011100111001101001011111101); #20
	MCMC_indirect_write(11'd1553, 68'b11001110010011000111001100111001011110100111011011011101110100110011); #20
	MCMC_indirect_write(11'd1554, 68'b11101101001001010111010011101100101101101010100010011011100100110101); #20
	MCMC_indirect_write(11'd1555, 68'b11111000000011011000000000000000010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1556, 68'b10100001000100001100111101101101001001001011010001110100101111110001); #20
	MCMC_indirect_write(11'd1557, 68'b10100011111101111100101101100101011000000110110100110001000001111001); #20
	MCMC_indirect_write(11'd1558, 68'b11101101100111110111101101110101011111001010011000011110111100111111); #20
	MCMC_indirect_write(11'd1559, 68'b11000001000101110100011000010000111010001010111010110110101001101000); #20
	MCMC_indirect_write(11'd1560, 68'b10110000111000111101010100011100001001000110010110110100011111000011); #20
	MCMC_indirect_write(11'd1561, 68'b10000000000000000100000000000000000100000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1562, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1563, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1564, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1565, 68'b01010100100000000010101100001100010100001100001111101010100100011001); #20
	MCMC_indirect_write(11'd1566, 68'b10000101110110111110000100110011111010001001010011010011001001110001); #20
	MCMC_indirect_write(11'd1567, 68'b01101000001010001100000100001010101000101111001100101000100011111111); #20
	MCMC_indirect_write(11'd1568, 68'b01001011101010010010101111001110100100010111100110000011000110011111); #20
	MCMC_indirect_write(11'd1569, 68'b10001011100010101100010010001011010111110111100111001001111001010110); #20
	MCMC_indirect_write(11'd1570, 68'b10110100100100011110010110011011011100100111100100110100001110000000); #20
	MCMC_indirect_write(11'd1571, 68'b10010101000101110011010101010000001000011101100110110001100101111111); #20
	MCMC_indirect_write(11'd1572, 68'b11100010000000011111001101100011111100101011010000111111010011011000); #20
	MCMC_indirect_write(11'd1573, 68'b11001100000101010101011100110000101011011001011100010110101000001111); #20
	MCMC_indirect_write(11'd1574, 68'b01110110100110001011111100111011111001111001100111110100010011110110); #20
	MCMC_indirect_write(11'd1575, 68'b11100000101111111111010000001000101111111100011101011110110011100000); #20
	MCMC_indirect_write(11'd1576, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1577, 68'b00001010010100001000101110101110000000100010010011100001010010000101); #20
	MCMC_indirect_write(11'd1578, 68'b10011001001110100101001001010101111011101110010011011011101100011101); #20
	MCMC_indirect_write(11'd1579, 68'b11001000111101100110010111011001011100001111111101110110011011110000); #20
	MCMC_indirect_write(11'd1580, 68'b11100100000111000110110000110111101100000011001110110110001100010001); #20
	MCMC_indirect_write(11'd1581, 68'b01110011110101011011110100001111000110110000001110110001111111011010); #20
	MCMC_indirect_write(11'd1582, 68'b10001000111010101100111100110111110111101000111001101111110010011011); #20
	MCMC_indirect_write(11'd1583, 68'b10000000000000000010000000000000000111111110100101011111111010011010); #20
	MCMC_indirect_write(11'd1584, 68'b01101101000000011011101111001111011001011110011001110111010100111111); #20
	MCMC_indirect_write(11'd1585, 68'b01110100011111101011100101010010010110000011100100001000011000110000); #20
	MCMC_indirect_write(11'd1586, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1587, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1588, 68'b11001010100010101101110110010000011000011001011010110010001010100111); #20
	MCMC_indirect_write(11'd1589, 68'b11111011111001001100000000000000000111110011011111011000000000000000); #20
	MCMC_indirect_write(11'd1590, 68'b10000000000000000010000000000000000100000000000000001000000000000000); #20
	MCMC_indirect_write(11'd1591, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1592, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1593, 68'b01110100010110001100001101110010011010100111111001010110011100101100); #20
	MCMC_indirect_write(11'd1594, 68'b11101001011111100100000000000000000100000000000000001111111110000010); #20
	MCMC_indirect_write(11'd1595, 68'b10000101000001111011011111010010110111011100101110101010110111101010); #20
	MCMC_indirect_write(11'd1596, 68'b11010111000100110110010110100100001101000101110000111000011100100111); #20
	MCMC_indirect_write(11'd1597, 68'b11000001110100010100011001100101011001110000110000001101111011010110); #20
	MCMC_indirect_write(11'd1598, 68'b10111100100001100110100111011001011101011001010000010111111110101010); #20
	MCMC_indirect_write(11'd1599, 68'b10000000000000000100000000000000001000000000000000011111100000011010); #20
	MCMC_indirect_write(11'd1600, 68'b11001000000000000110010000000000001100100000000000011001000000000000); #20
	MCMC_indirect_write(11'd1601, 68'b11011010111011110110110000001101011101000010101000111001111110011100); #20
	MCMC_indirect_write(11'd1602, 68'b11001111001110011110101001001001101011011111111101011011010010110011); #20
	MCMC_indirect_write(11'd1603, 68'b11100011001001011110010000111000101110011111000110111100011111100110); #20
	MCMC_indirect_write(11'd1604, 68'b10101100111000010101111110001011011110001100110000111000001111001011); #20
	MCMC_indirect_write(11'd1605, 68'b10101001110110000111001010000010001111101001010111011100001000110010); #20
	MCMC_indirect_write(11'd1606, 68'b10001101110111111100110010101111101010110001100001011000010000110111); #20
	MCMC_indirect_write(11'd1607, 68'b11011010111000110110000011000001001100110001010001011011011110000010); #20
	MCMC_indirect_write(11'd1608, 68'b10101011100100100101001000000010001001100100110111010001101100101101); #20
	MCMC_indirect_write(11'd1609, 68'b10110110101111000110101111100110111101101100100101111001011110001010); #20
	MCMC_indirect_write(11'd1610, 68'b11011101001101100111011100011010111101101100010101111010011010110101); #20
	MCMC_indirect_write(11'd1611, 68'b10100010010110111101010111011111110111001100111011001100011010000100); #20
	MCMC_indirect_write(11'd1612, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1613, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1614, 68'b01101010011001110011100011001010000100111101111110001000010010011001); #20
	MCMC_indirect_write(11'd1615, 68'b11001101000000111101001101100011011100011010101100110100101000001000); #20
	MCMC_indirect_write(11'd1616, 68'b11010110100111110110100010110000011101111000010001011011100001111110); #20
	MCMC_indirect_write(11'd1617, 68'b10000010100110101100110011001111111001011000101010010011010010111011); #20
	MCMC_indirect_write(11'd1618, 68'b11100000011010011110100001110101001010111000110000110010011110101110); #20
	MCMC_indirect_write(11'd1619, 68'b10110001101100000111001011000010001111010100000001111001111100010111); #20
	MCMC_indirect_write(11'd1620, 68'b01101001010111101010101111010101100100011011100010101010010010111100); #20
	MCMC_indirect_write(11'd1621, 68'b11010010100111001111101101101101101111001001111110011011110100000001); #20
	MCMC_indirect_write(11'd1622, 68'b10111101100011000101111001111011101100100100000000110101111111111100); #20
	MCMC_indirect_write(11'd1623, 68'b10111110100111110100010000001111011001011000000101101110010110000011); #20
	MCMC_indirect_write(11'd1624, 68'b10010100111000000101001001000001111000111000000111010100111001001010); #20
	MCMC_indirect_write(11'd1625, 68'b10000000000000000011101101001000110110000101000111111111101001110011); #20
	MCMC_indirect_write(11'd1626, 68'b11101000011100001111000010101100001111111010101101110000000000000000); #20
	MCMC_indirect_write(11'd1627, 68'b11110010001001111000000000000000010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1628, 68'b10000000000000001000000000000000010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1629, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1630, 68'b11110001111100100111101011110010011111101101000110011111111011111001); #20
	MCMC_indirect_write(11'd1631, 68'b11101010010000010111010011100011001000000000000000001101010011100100); #20
	MCMC_indirect_write(11'd1632, 68'b11001010110101001101110110000111101011100100100010011010101001100100); #20
	MCMC_indirect_write(11'd1633, 68'b10111110011111110101111001111101011011001101001100110100011000000000); #20
	MCMC_indirect_write(11'd1634, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1635, 68'b10111001111001101110001011111101001100110101001110111110001110011101); #20
	MCMC_indirect_write(11'd1636, 68'b01001010000101000011101001011011011000001100110000110000010011100110); #20
	MCMC_indirect_write(11'd1637, 68'b00000000000000000000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1638, 68'b10100001001010110100001010100100001001010101101011110100111010010011); #20
	MCMC_indirect_write(11'd1639, 68'b10111110100100111101011101110110001010000001010010010010011001100001); #20
	MCMC_indirect_write(11'd1640, 68'b10000000000000000111100100001101110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1641, 68'b10110110110100000110110010101100011101101001011101110111110000110101); #20
	MCMC_indirect_write(11'd1642, 68'b10111000011111111101000100011101011100010101111100010101111010001111); #20
	MCMC_indirect_write(11'd1643, 68'b11100000001100100110010110111000101110011010000101111011100110101011); #20
	MCMC_indirect_write(11'd1644, 68'b10000000000000000100000000000000001000000000000000011101001110010011); #20
	MCMC_indirect_write(11'd1645, 68'b01100000110110100001100101100110010000010101100111000010110011100111); #20
	MCMC_indirect_write(11'd1646, 68'b11010111100001100101010010111010101010000100100110001110000101101010); #20
	MCMC_indirect_write(11'd1647, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1648, 68'b01100110101010110010111100001101000110101010111110001010101100001001); #20
	MCMC_indirect_write(11'd1649, 68'b01110010111011101010111101110010110110001000101011001010101101000010); #20
	MCMC_indirect_write(11'd1650, 68'b10101000101101110110001010001000001000000000000000011011010101111010); #20
	MCMC_indirect_write(11'd1651, 68'b11001010011000111101101101110111101000110011010011110010011110110001); #20
	MCMC_indirect_write(11'd1652, 68'b10101011110100010110001001011110001011011110111010011001100100110101); #20
	MCMC_indirect_write(11'd1653, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1654, 68'b11111101101010100111010000010101101000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1655, 68'b00011110000000101001110000100101100010110000101010100001001010001010); #20
	MCMC_indirect_write(11'd1656, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1657, 68'b11100101110100001110011111110010101110010000101000011100011110100011); #20
	MCMC_indirect_write(11'd1658, 68'b11101100101011110110101110000010001100110011101001111111100111111010); #20
	MCMC_indirect_write(11'd1659, 68'b10100101101111100101100000101001111100101100000100111010110011011011); #20
	MCMC_indirect_write(11'd1660, 68'b10000000000000000100000000000000001000000000000000011111110111100100); #20
	MCMC_indirect_write(11'd1661, 68'b10110010010100010110000000100010111101111001100111011100010000011101); #20
	MCMC_indirect_write(11'd1662, 68'b10001110001101001011011110111101110111010011110001101111110101010111); #20
	MCMC_indirect_write(11'd1663, 68'b10000000000000000111010100111110001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1664, 68'b11010000000000000110100000000000001101000000000000011010000000000000); #20
	MCMC_indirect_write(11'd1665, 68'b11001011000001000110011100100111111011111110010011111001100010101001); #20
	MCMC_indirect_write(11'd1666, 68'b11010010000100100111001010100001111101100101111100011011110100010010); #20
	MCMC_indirect_write(11'd1667, 68'b11011010111110110111000010010010001101011011001110111000100100100010); #20
	MCMC_indirect_write(11'd1668, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1669, 68'b11010110011101011110011100100001101000000000000000011111010100101011); #20
	MCMC_indirect_write(11'd1670, 68'b11011100100010110110010010000100101110010101111011011100010001100110); #20
	MCMC_indirect_write(11'd1671, 68'b11010101011001111111000111101111111110100101111101011111110111101100); #20
	MCMC_indirect_write(11'd1672, 68'b11111011000101001110111111001010110000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1673, 68'b11011110110000011111111111100011111000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1674, 68'b11101000000111110110011000110000101110111001100011111010011111111101); #20
	MCMC_indirect_write(11'd1675, 68'b01100001100110001011000011111011101000011100001001110111000100111111); #20
	MCMC_indirect_write(11'd1676, 68'b11000100100010001111000101010000011011100011101100010110111111010100); #20
	MCMC_indirect_write(11'd1677, 68'b01100100111110000011011111011011100101010111000011001101001010100000); #20
	MCMC_indirect_write(11'd1678, 68'b10101011110001011100001110101101011001000001111000110001001011101110); #20
	MCMC_indirect_write(11'd1679, 68'b10111011111011100100100111001101011010001000010000010101010111100100); #20
	MCMC_indirect_write(11'd1680, 68'b11101001010110011110111011010100101111100101100010111101111010111111); #20
	MCMC_indirect_write(11'd1681, 68'b11100010100110101110010000110101001010110111111001010001100000111111); #20
	MCMC_indirect_write(11'd1682, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1683, 68'b11110001101111001110101111000000011101001000010101010011111000101010); #20
	MCMC_indirect_write(11'd1684, 68'b11110011100001011111010011111111011111100111000011111110010000010101); #20
	MCMC_indirect_write(11'd1685, 68'b10000000000000000100000000000000001110111101010110111000010100111110); #20
	MCMC_indirect_write(11'd1686, 68'b01010101111101110011001010010110010100111111100011000110010100111000); #20
	MCMC_indirect_write(11'd1687, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1688, 68'b11010110001100111100000000000000001110010000101100011010100001000101); #20
	MCMC_indirect_write(11'd1689, 68'b00010101010110110000000000000000000000000000000000000000000000000000); #20
	MCMC_indirect_write(11'd1690, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1691, 68'b11111010010001110100000000000000001111111100100010010000000000000000); #20
	MCMC_indirect_write(11'd1692, 68'b10001010011011010011111101010110100100110010000010100111100111010111); #20
	MCMC_indirect_write(11'd1693, 68'b01100001100111000010110011001001110110001010101101101010010110000010); #20
	MCMC_indirect_write(11'd1694, 68'b01011011111100000010001000010100010100111011111011001010100110100000); #20
	MCMC_indirect_write(11'd1695, 68'b11001100101011100101101001110001101100001011111000110010110001000101); #20
	MCMC_indirect_write(11'd1696, 68'b10010100111110011101010001010000101000101000010110110011010110111100); #20
	MCMC_indirect_write(11'd1697, 68'b01100101001100000011110101101100101000101101000111010001010100000010); #20
	MCMC_indirect_write(11'd1698, 68'b10110001011000100110010000110110111101001001010100110010111101100010); #20
	MCMC_indirect_write(11'd1699, 68'b11110100110001101111111010101000001111111110111110011110100110010000); #20
	MCMC_indirect_write(11'd1700, 68'b00011000001001011000110000101111000000000000000000000010001110011101); #20
	MCMC_indirect_write(11'd1701, 68'b11000110111000011110001100011110101100101110001110111011111001001111); #20
	MCMC_indirect_write(11'd1702, 68'b11110111010011101100000000000000001000000000000000011111010100100010); #20
	MCMC_indirect_write(11'd1703, 68'b10100001010111011100101110100011001000110100101001001101001110100111); #20
	MCMC_indirect_write(11'd1704, 68'b10011000010111101101001100000000111011000001101011011011110100011000); #20
	MCMC_indirect_write(11'd1705, 68'b10001100010110000100001110111010011000001011001101010011111100010100); #20
	MCMC_indirect_write(11'd1706, 68'b01110100100011100100001000010001100111010111010000101111101100110001); #20
	MCMC_indirect_write(11'd1707, 68'b11010010001110111111101101000001011111011111101110100000000000000000); #20
	MCMC_indirect_write(11'd1708, 68'b11100011000000111111010001011010101110011100110110110000000000000000); #20
	MCMC_indirect_write(11'd1709, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1710, 68'b10010010001000100100110101110110001000110010101011110001110011000100); #20
	MCMC_indirect_write(11'd1711, 68'b10101111010010111011110111010111100110110011100100001000100001001110); #20
	MCMC_indirect_write(11'd1712, 68'b11010110110011011110100001001001001101000001010101111001101011001100); #20
	MCMC_indirect_write(11'd1713, 68'b10110111101000101100000110111000110110110101110000101011110101101110); #20
	MCMC_indirect_write(11'd1714, 68'b01110000010000111011100111011000010100011101010001100100111101101010); #20
	MCMC_indirect_write(11'd1715, 68'b01000011101000100001000011101101010011100000110011001000010110111011); #20
	MCMC_indirect_write(11'd1716, 68'b11010101011111101110111100110110101101110010010100111000110001100111); #20
	MCMC_indirect_write(11'd1717, 68'b10010000001100101101000101111011101010100000100101110100010010111101); #20
	MCMC_indirect_write(11'd1718, 68'b11011000001110001110010011110100101011001101001010011011111011110111); #20
	MCMC_indirect_write(11'd1719, 68'b11011111110000001101110001110101001011010010101001010111100011101111); #20
	MCMC_indirect_write(11'd1720, 68'b11100110101011000111101001010111101111010101100001011101010101111001); #20
	MCMC_indirect_write(11'd1721, 68'b11011110100100011100110101110001111110011010111000100000000000000000); #20
	MCMC_indirect_write(11'd1722, 68'b11100010100111100111010101001110011000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1723, 68'b01110011100111110011011000011010111001010001100001011001111001010011); #20
	MCMC_indirect_write(11'd1724, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1725, 68'b01011000101011001011110110010111110111001100111110110000111101100010); #20
	MCMC_indirect_write(11'd1726, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1727, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1728, 68'b11011000000000000110110000000000001101100000000000011011000000000000); #20
	MCMC_indirect_write(11'd1729, 68'b11010100100001010110000010110011011101111101100100011010001010011011); #20
	MCMC_indirect_write(11'd1730, 68'b11001100110010111111010101000111111100111000111000111011111010010110); #20
	MCMC_indirect_write(11'd1731, 68'b11101111011001000110111010011011111101101010010111111111001010001001); #20
	MCMC_indirect_write(11'd1732, 68'b11011101001010001110101101010100001110101110011110111001101000011000); #20
	MCMC_indirect_write(11'd1733, 68'b10000000000000000100000000000000001110111011011111011110101110110110); #20
	MCMC_indirect_write(11'd1734, 68'b10101010110101001101110000001000111011011010011010011010101001100110); #20
	MCMC_indirect_write(11'd1735, 68'b10111101111011010110100001101101011101000001011011010100010111101000); #20
	MCMC_indirect_write(11'd1736, 68'b11100011011110100111011100001110011000000000000000011111101011101100); #20
	MCMC_indirect_write(11'd1737, 68'b00011111000101010000100010110011000000000100011110000000000000000000); #20
	MCMC_indirect_write(11'd1738, 68'b11000000000011001110000001111100001100111011101010011000110101111001); #20
	MCMC_indirect_write(11'd1739, 68'b11110010110101110111110111010001011110010101001111011100111100111100); #20
	MCMC_indirect_write(11'd1740, 68'b11101100001101110111011111001110011110000011101110111100110011111111); #20
	MCMC_indirect_write(11'd1741, 68'b11110011111110011110010000010101001110010011010110111101001011111101); #20
	MCMC_indirect_write(11'd1742, 68'b10110001001100111101011010100010011100111000000100111011000111011111); #20
	MCMC_indirect_write(11'd1743, 68'b11101001111011011111011000111110011110101111001011111011111001111000); #20
	MCMC_indirect_write(11'd1744, 68'b01101110011011010011011010101010100110011110111010001111110100000100); #20
	MCMC_indirect_write(11'd1745, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1746, 68'b11000011110111101101110000110000001000101111011100001111111010011111); #20
	MCMC_indirect_write(11'd1747, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1748, 68'b11110100010011110101111110101011111101111011110111111110000000100011); #20
	MCMC_indirect_write(11'd1749, 68'b10001111101111100101000010010000010111010011001011101110001000011111); #20
	MCMC_indirect_write(11'd1750, 68'b10100000000111100100110011000011001011000101011111011001000000011111); #20
	MCMC_indirect_write(11'd1751, 68'b11100011110110000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1752, 68'b11010010111011100101111011001010101010100101110000110001000000111010); #20
	MCMC_indirect_write(11'd1753, 68'b10000000000000000100000000000000001111101101001101010000000000000000); #20
	MCMC_indirect_write(11'd1754, 68'b11011001010001011111011110100000011111110101111101011101001011111110); #20
	MCMC_indirect_write(11'd1755, 68'b11011100110011100111101101101101111111101001010000110000000000000000); #20
	MCMC_indirect_write(11'd1756, 68'b10000000111111001100111000011010001000010011000100001100011110001010); #20
	MCMC_indirect_write(11'd1757, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1758, 68'b11101011101100001110010010010101101100101010101100110110101101001110); #20
	MCMC_indirect_write(11'd1759, 68'b10101010011100110101011001000110011010001111100100101111111011011110); #20
	MCMC_indirect_write(11'd1760, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1761, 68'b10010001011000101100111011110001001100011010010000011010101101001111); #20
	MCMC_indirect_write(11'd1762, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1763, 68'b00100101010011101001100001100110000010011001001101100001101100000111); #20
	MCMC_indirect_write(11'd1764, 68'b11000111001100011111000110010001001111101100011101111000000001100101); #20
	MCMC_indirect_write(11'd1765, 68'b01100011101000000100101111001101001000011110010000110001011101010101); #20
	MCMC_indirect_write(11'd1766, 68'b11000100011011011111010111101111011100110101010000011010110011111110); #20
	MCMC_indirect_write(11'd1767, 68'b11010100011001001100100101111110111110111100000011100000000000000000); #20
	MCMC_indirect_write(11'd1768, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1769, 68'b11101001011000011000000000000000010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1770, 68'b10001100001111100101101110100111111011111000110000110101111011000010); #20
	MCMC_indirect_write(11'd1771, 68'b10100101001000101101110110000110111110001001101101011110000011000101); #20
	MCMC_indirect_write(11'd1772, 68'b11010001001001001110110101010111001110111110110111111010111111011110); #20
	MCMC_indirect_write(11'd1773, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1774, 68'b10010101100100110011111010011111000110000011100111101110001100100101); #20
	MCMC_indirect_write(11'd1775, 68'b10100110111011010101011011001111101100100000101011011010000010101000); #20
	MCMC_indirect_write(11'd1776, 68'b10000111000011011010111101011000010111111010001100101011000100100011); #20
	MCMC_indirect_write(11'd1777, 68'b10000000000000000010000000000000000111000100010010110000000000000000); #20
	MCMC_indirect_write(11'd1778, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1779, 68'b01111110000010100011101010101001110110001001111111100111000100000011); #20
	MCMC_indirect_write(11'd1780, 68'b10101100000101010101001101001101111000111110100110110010111001000011); #20
	MCMC_indirect_write(11'd1781, 68'b11110110111001101111100111011100001110101010110101111010001111101100); #20
	MCMC_indirect_write(11'd1782, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1783, 68'b10110000011000111100100011111100001000110010111011110001100110110100); #20
	MCMC_indirect_write(11'd1784, 68'b00101001010010100010000010000101010100011011100100001101011101000001); #20
	MCMC_indirect_write(11'd1785, 68'b11110100101100100110101011011111011111111111111111110000000000000000); #20
	MCMC_indirect_write(11'd1786, 68'b11000001111010110110011011100100001100010010100100110110100010011000); #20
	MCMC_indirect_write(11'd1787, 68'b11110101100011011111100011001011101110110101001000111100111011110011); #20
	MCMC_indirect_write(11'd1788, 68'b10000111110110001101101111111000011010101011110001010101100010111010); #20
	MCMC_indirect_write(11'd1789, 68'b10001101001110000100000010101011101000111011110000110001001100110111); #20
	MCMC_indirect_write(11'd1790, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1791, 68'b11011111100010101100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1792, 68'b11100000000000000111000000000000001110000000000000011100000000000000); #20
	MCMC_indirect_write(11'd1793, 68'b11011100111010010110111000000001111110101011000111111100101100100011); #20
	MCMC_indirect_write(11'd1794, 68'b11011000111010001111010000110101111111100011111101111101011000110010); #20
	MCMC_indirect_write(11'd1795, 68'b11011001101000111111000010101011011111001101100110011111110010000011); #20
	MCMC_indirect_write(11'd1796, 68'b10000000000000000010000000000000000111101001110111011110111110000010); #20
	MCMC_indirect_write(11'd1797, 68'b11111100100001111111010011101000011000000000000000011111111001111001); #20
	MCMC_indirect_write(11'd1798, 68'b11001101110110001110001010111101111100111101001011011010001110001000); #20
	MCMC_indirect_write(11'd1799, 68'b11100001000001101111011010101100101110011111100110111010110010000110); #20
	MCMC_indirect_write(11'd1800, 68'b10000000000000000100000000000000001110101101110011111010000110010011); #20
	MCMC_indirect_write(11'd1801, 68'b11101101000101100111000000111111001100111111010110011001011011011011); #20
	MCMC_indirect_write(11'd1802, 68'b11001111110010011110100111110001011101101111011001111100110000111011); #20
	MCMC_indirect_write(11'd1803, 68'b11101101111100100111001100000010111101010011101000111110101011110111); #20
	MCMC_indirect_write(11'd1804, 68'b11011110111110101110000111011111011101101000011101111011001101110010); #20
	MCMC_indirect_write(11'd1805, 68'b11100110100001111110110101001111001100110010101100011100010011100111); #20
	MCMC_indirect_write(11'd1806, 68'b11001101111110010110010001101011001101111110011111110110110110011001); #20
	MCMC_indirect_write(11'd1807, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1808, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1809, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1810, 68'b10000100010001101100011111111011111001110001110100110010100111011100); #20
	MCMC_indirect_write(11'd1811, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1812, 68'b11000000110001110100100001001110111010010111101010010101101001110011); #20
	MCMC_indirect_write(11'd1813, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1814, 68'b11110011100101010110011100100111101011000000101011010110000001110101); #20
	MCMC_indirect_write(11'd1815, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1816, 68'b10010010000011111101011100011100011001011100011011011010001011000110); #20
	MCMC_indirect_write(11'd1817, 68'b11100101100111100111001110011001011110101100110001011011011000010001); #20
	MCMC_indirect_write(11'd1818, 68'b10100111001101001101100101011001101100011001101111110111100001111000); #20
	MCMC_indirect_write(11'd1819, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1820, 68'b11100010010100110110101000000101111100100111010100010100101001001000); #20
	MCMC_indirect_write(11'd1821, 68'b10111001110000110100011100000101111000100000001110001101111011100111); #20
	MCMC_indirect_write(11'd1822, 68'b01111000111011101011101011100001101001110011110100110100010010001110); #20
	MCMC_indirect_write(11'd1823, 68'b10001001011011100011010011110110100111001101001100110000010110000010); #20
	MCMC_indirect_write(11'd1824, 68'b11001110110111101101111100110001111011111111001001010110000011110000); #20
	MCMC_indirect_write(11'd1825, 68'b10011000100011100101011110010001011001011110000100101110101001100100); #20
	MCMC_indirect_write(11'd1826, 68'b11001100111101111101110001111100011100001100101101010010000010110100); #20
	MCMC_indirect_write(11'd1827, 68'b01100101101101100011100000100110110101101000011001110000010110110010); #20
	MCMC_indirect_write(11'd1828, 68'b10110001001101111101100101001101001010110110000011010010000110010110); #20
	MCMC_indirect_write(11'd1829, 68'b10011001000101000101110110001001101011100100011100111110001101100000); #20
	MCMC_indirect_write(11'd1830, 68'b10000000000000000100000000000000001101110111111010010111101110000001); #20
	MCMC_indirect_write(11'd1831, 68'b10010111001111100100100100110111001001110011010011001111100100101101); #20
	MCMC_indirect_write(11'd1832, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1833, 68'b10100111010101001101100000000010101001110000111011110001001110011100); #20
	MCMC_indirect_write(11'd1834, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1835, 68'b01100010110000101010101001011111000101100010110011010000100110111011); #20
	MCMC_indirect_write(11'd1836, 68'b11011101010100110111011101011110011111100001111000011110001000001011); #20
	MCMC_indirect_write(11'd1837, 68'b11011010110000000110011111100110111100111110001001110000000000000000); #20
	MCMC_indirect_write(11'd1838, 68'b10010101001111100101100011000000011010001011100111010011111101010011); #20
	MCMC_indirect_write(11'd1839, 68'b11001111111111010111100010000110001111001101111110010000000000000000); #20
	MCMC_indirect_write(11'd1840, 68'b11010001111110111111100110111101101110100100110100110000000000000000); #20
	MCMC_indirect_write(11'd1841, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1842, 68'b10000000000000000111101011000000111111011111110001011111000011000101); #20
	MCMC_indirect_write(11'd1843, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1844, 68'b11111010100111000110111111000011011111101111010100110000000000000000); #20
	MCMC_indirect_write(11'd1845, 68'b10000000000000000111110001000001111111010011100101011001111111111100); #20
	MCMC_indirect_write(11'd1846, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1847, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1848, 68'b11110101011110101100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1849, 68'b11111011110101111100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1850, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1851, 68'b11010010000101011111001011101101101110001101011010111101001011011001); #20
	MCMC_indirect_write(11'd1852, 68'b01000111110000100010010111111001010010111101100001101010010011110100); #20
	MCMC_indirect_write(11'd1853, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1854, 68'b10000000000000000100000000000000001000000000000000011110101111101010); #20
	MCMC_indirect_write(11'd1855, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1856, 68'b11101000000000000111010000000000001110100000000000011101000000000000); #20
	MCMC_indirect_write(11'd1857, 68'b11100111100000110111001001100110001110000100010111011101111001000011); #20
	MCMC_indirect_write(11'd1858, 68'b11101001111000001111010000110101011110111101000000111111011110011101); #20
	MCMC_indirect_write(11'd1859, 68'b10111100111100100110000010011100011110101110110111010110111000100110); #20
	MCMC_indirect_write(11'd1860, 68'b11101001000011101110110111110001001011110110111011010111110110001000); #20
	MCMC_indirect_write(11'd1861, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1862, 68'b11110000110000111000000000000000010000000000000000011111011001001011); #20
	MCMC_indirect_write(11'd1863, 68'b10000000000000000100000000000000000100000000000000011110000011110011); #20
	MCMC_indirect_write(11'd1864, 68'b10000000000000000010000000000000000111111100010111111111001011010110); #20
	MCMC_indirect_write(11'd1865, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1866, 68'b11010110010001101111010011001111111100010010010110011101110111000011); #20
	MCMC_indirect_write(11'd1867, 68'b10110010000110101100110001100110101010001000111101010111111101101001); #20
	MCMC_indirect_write(11'd1868, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1869, 68'b10000000000000000111110110101111111111011010100011011111010001101100); #20
	MCMC_indirect_write(11'd1870, 68'b11010101100001101110110101110010111101110110000001100000000000000000); #20
	MCMC_indirect_write(11'd1871, 68'b11111000010001111111001111110101111110100110001001111111001001101111); #20
	MCMC_indirect_write(11'd1872, 68'b11110001101101001100000000000000001000000000000000011110001111010100); #20
	MCMC_indirect_write(11'd1873, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1874, 68'b11101111110011011111011111101001010000000000000000100000000000000000); #20
	MCMC_indirect_write(11'd1875, 68'b11010000101010000101100110100111011011000001110110010101011001011010); #20
	MCMC_indirect_write(11'd1876, 68'b11001001000011010101101000011100001000001100010110001110000010100110); #20
	MCMC_indirect_write(11'd1877, 68'b11011110000100001110010000011001111011111000010011110011001111001010); #20
	MCMC_indirect_write(11'd1878, 68'b01011001001100101001011111100110110101111000110100001101111111001101); #20
	MCMC_indirect_write(11'd1879, 68'b11101010100100001101110000000010010111000110010110001111011101011100); #20
	MCMC_indirect_write(11'd1880, 68'b10111010101011010100100110010001111100110100011111010111100101001010); #20
	MCMC_indirect_write(11'd1881, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1882, 68'b10000000000000000111010010111110001111110010010001011111011110000001); #20
	MCMC_indirect_write(11'd1883, 68'b11110110101001001111010010101100001111010101111010111111111011110010); #20
	MCMC_indirect_write(11'd1884, 68'b10011101110001111110001111111010101100110100100101111100001010010001); #20
	MCMC_indirect_write(11'd1885, 68'b10011101011010010101001011011001001010111001001011111001100110011010); #20
	MCMC_indirect_write(11'd1886, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1887, 68'b10000000000000000100000000000000001111111011000111011110101111001101); #20
	MCMC_indirect_write(11'd1888, 68'b10101000100010100101111111010001001011111100000110011010001001011101); #20
	MCMC_indirect_write(11'd1889, 68'b11111100000011101111110011011000110000000000000000011101110000100111); #20
	MCMC_indirect_write(11'd1890, 68'b11100001100001110111001000110110011101111001011000110101010100110010); #20
	MCMC_indirect_write(11'd1891, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1892, 68'b11101111100000110100000000000000001111111101111000010000000000000000); #20
	MCMC_indirect_write(11'd1893, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1894, 68'b10011101010011111100100101111000011101001101111111110100001000100101); #20
	MCMC_indirect_write(11'd1895, 68'b11010000001011110110101000011001111100110011000011010110110110101100); #20
	MCMC_indirect_write(11'd1896, 68'b10010010101110010100011010001111011000110110001001010000100000011001); #20
	MCMC_indirect_write(11'd1897, 68'b11110111000110111111001010000000011111010001000000110000000000000000); #20
	MCMC_indirect_write(11'd1898, 68'b11010011000010011101010000111110111110001010101001100000000000000000); #20
	MCMC_indirect_write(11'd1899, 68'b10000000000000000011100001011101101111100011110110010000000000000000); #20
	MCMC_indirect_write(11'd1900, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1901, 68'b10110000101011000101111011101000001100100010110000011001111110001000); #20
	MCMC_indirect_write(11'd1902, 68'b10100011101001100100110101101011111011010011011111110110010010101010); #20
	MCMC_indirect_write(11'd1903, 68'b10100100010111110101001011101010111010100111111100010110100110110001); #20
	MCMC_indirect_write(11'd1904, 68'b11101001011111010111000010100100011110111100100110011010011111001110); #20
	MCMC_indirect_write(11'd1905, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1906, 68'b01110010101011010100000100100110101001001101111000110110110111000100); #20
	MCMC_indirect_write(11'd1907, 68'b11000111000101000110111010011011101101100010011100110111100100001001); #20
	MCMC_indirect_write(11'd1908, 68'b11010000110001010111010010111100101011010100101111010101111100011100); #20
	MCMC_indirect_write(11'd1909, 68'b11111000010011101110111010000000011111100011101001011011100100101111); #20
	MCMC_indirect_write(11'd1910, 68'b11101000011110101111110011100100001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1911, 68'b11110010101111000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1912, 68'b11010010110101000111010101001110011101111010100111010101101011110000); #20
	MCMC_indirect_write(11'd1913, 68'b01001010011010010010011001110110110011001111011011000110101111101011); #20
	MCMC_indirect_write(11'd1914, 68'b10000000000000000100000000000000001000000000000000011111000001100100); #20
	MCMC_indirect_write(11'd1915, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1916, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1917, 68'b11110111011000011100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1918, 68'b11011011110100100110010001111010111100001010101000111000000001110010); #20
	MCMC_indirect_write(11'd1919, 68'b10000000000000000100000000000000001111100010001100011100101111101010); #20
	MCMC_indirect_write(11'd1920, 68'b11110000000000000111100000000000001111000000000000011110000000000000); #20
	MCMC_indirect_write(11'd1921, 68'b11101100101110110111100110010011101111001001010000011101111001100111); #20
	MCMC_indirect_write(11'd1922, 68'b11101110000001011111101011101010001110111010011101111111010010110001); #20
	MCMC_indirect_write(11'd1923, 68'b10000000000000000100000000000000001000000000000000011100101011010110); #20
	MCMC_indirect_write(11'd1924, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1925, 68'b11100011101100010111111010101100011000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1926, 68'b11110111110111001100000000000000001111000110101101011101011011111000); #20
	MCMC_indirect_write(11'd1927, 68'b11001000000011101110011100110111111101110101010000111011101111110000); #20
	MCMC_indirect_write(11'd1928, 68'b10101001001010011110100011001100011001110111111100010100011011101001); #20
	MCMC_indirect_write(11'd1929, 68'b10111010000101100111010011011100011110101100101000011110100010101110); #20
	MCMC_indirect_write(11'd1930, 68'b10111111100000010110001001001011101101011010101100111100111000011111); #20
	MCMC_indirect_write(11'd1931, 68'b11110101001100010111101100011001011110101000010111111000101111011011); #20
	MCMC_indirect_write(11'd1932, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1933, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1934, 68'b11101111010001011000000000000000011111000111010111100000000000000000); #20
	MCMC_indirect_write(11'd1935, 68'b01100011011010000011111011010000110111010101101000010001001111100010); #20
	MCMC_indirect_write(11'd1936, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1937, 68'b11010101110110011111000101001111001110110111011010111011011111010001); #20
	MCMC_indirect_write(11'd1938, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1939, 68'b11001001001001001101010000110111111001001101101101010001110110101101); #20
	MCMC_indirect_write(11'd1940, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1941, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1942, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1943, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1944, 68'b11010000000000100110100101111111001100101001001101011010101100110000); #20
	MCMC_indirect_write(11'd1945, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1946, 68'b11100111001110010100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1947, 68'b11100111111011101111000100110101101101000001000101010101101111111010); #20
	MCMC_indirect_write(11'd1948, 68'b11001110100000001111011101101100001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1949, 68'b11010010010000001110100011000010001101010001010101011010011001010101); #20
	MCMC_indirect_write(11'd1950, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1951, 68'b10001111101001001100100000100001010110101101010110101010110100100100); #20
	MCMC_indirect_write(11'd1952, 68'b10101110011101101101111101101011011010111000111101010111101101111110); #20
	MCMC_indirect_write(11'd1953, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1954, 68'b10010011101001011100011111111111011010110000000111111001001011010001); #20
	MCMC_indirect_write(11'd1955, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1956, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1957, 68'b11111100001001111111001100100010011100100110110110110011110101000100); #20
	MCMC_indirect_write(11'd1958, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1959, 68'b11110111100011000111001010011001001111000011100101111110011010110001); #20
	MCMC_indirect_write(11'd1960, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1961, 68'b10001001011010011011101101110100101000110111000010110111000111101111); #20
	MCMC_indirect_write(11'd1962, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1963, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1964, 68'b10110011001001011101111001001001111011101011101100111101110100010011); #20
	MCMC_indirect_write(11'd1965, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1966, 68'b11000111100101110101001111001000011010101101000000110110011110100000); #20
	MCMC_indirect_write(11'd1967, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1968, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1969, 68'b00111101101100100010001110011110010001000010111011100010101001001111); #20
	MCMC_indirect_write(11'd1970, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1971, 68'b10000000000000000100000000000000001000000000000000011111110001111000); #20
	MCMC_indirect_write(11'd1972, 68'b11100101010010110100000000000000001110101111100110111100111011000100); #20
	MCMC_indirect_write(11'd1973, 68'b10000000000000000100000000000000001000000000000000011110001101011011); #20
	MCMC_indirect_write(11'd1974, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1975, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1976, 68'b01100110000010000011101010110010001000101000110000010001100101010000); #20
	MCMC_indirect_write(11'd1977, 68'b11110111000111110100000000000000001000000000000000010110000110110111); #20
	MCMC_indirect_write(11'd1978, 68'b10101101100100110101010110010000111010000010110011110100110110100010); #20
	MCMC_indirect_write(11'd1979, 68'b10011100110100011101110011000110011101001010111010111010101101010111); #20
	MCMC_indirect_write(11'd1980, 68'b10000000000000000100000000000000001110010110100101011111011011100000); #20
	MCMC_indirect_write(11'd1981, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1982, 68'b11100111001001101111110110010111001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1983, 68'b11011010100000010101111110001101111100011001001101010101010101101110); #20
	MCMC_indirect_write(11'd1984, 68'b11111000000000000111110000000000001111100000000000011111000000000000); #20
	MCMC_indirect_write(11'd1985, 68'b11111111110010010111100110000100111111111100110101110000000000000000); #20
	MCMC_indirect_write(11'd1986, 68'b11100001011010100111100101111101101110110000110010011101110100111000); #20
	MCMC_indirect_write(11'd1987, 68'b11100000110101001111111101011110111101001101011100111010100111011010); #20
	MCMC_indirect_write(11'd1988, 68'b11110111111011011111110101101100001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1989, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1990, 68'b11010110010100101100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1991, 68'b01111010111100001011011111010010010111010010001100001011100010000100); #20
	MCMC_indirect_write(11'd1992, 68'b11110010110000111111100111001110001110011111111000011110101011010000); #20
	MCMC_indirect_write(11'd1993, 68'b10011111000100110110000110011101101100000011100100010100010110001011); #20
	MCMC_indirect_write(11'd1994, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1995, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1996, 68'b11110000011101101100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd1997, 68'b10001111011100010100001000011011101010000100101101010010111001011001); #20
	MCMC_indirect_write(11'd1998, 68'b10010101101111111011111010111001001001110110101101001111001110110101); #20
	MCMC_indirect_write(11'd1999, 68'b11110110101110001110110111011110101110010010110110111100010101111100); #20
	MCMC_indirect_write(11'd2000, 68'b10000000000000000100000000000000001111000110110101011111101101001101); #20
	MCMC_indirect_write(11'd2001, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2002, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2003, 68'b11101101011110101110101001000011111100100100011111010010001100101100); #20
	MCMC_indirect_write(11'd2004, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2005, 68'b11010011111110101110101001001010111110001000100010011110000101100010); #20
	MCMC_indirect_write(11'd2006, 68'b11110010000111001100000000000000001000000000000000001110110111010101); #20
	MCMC_indirect_write(11'd2007, 68'b10010011010110111011011000001011101001101000000010001110110111111000); #20
	MCMC_indirect_write(11'd2008, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2009, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2010, 68'b11111111110001111100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2011, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2012, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2013, 68'b11010000101100010110101011011101011110100000110001111000110010111001); #20
	MCMC_indirect_write(11'd2014, 68'b10000000000000000100000000000000001000000000000000011100001111011011); #20
	MCMC_indirect_write(11'd2015, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2016, 68'b11111101010001010100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2017, 68'b01111000010100111100111010010001101001000011011101101111110110011001); #20
	MCMC_indirect_write(11'd2018, 68'b11010001011100011101110111111110111110010100100110111111010100100100); #20
	MCMC_indirect_write(11'd2019, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2020, 68'b10110111011111001101110110100001101001110011100100110010000110001011); #20
	MCMC_indirect_write(11'd2021, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2022, 68'b11011011011010101110001101000110101010010110110110010101011010111101); #20
	MCMC_indirect_write(11'd2023, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2024, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2025, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2026, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2027, 68'b11011100000101100111000000111100101101001100110101010111010110011011); #20
	MCMC_indirect_write(11'd2028, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2029, 68'b11110010100000001111001001101010111000000000000000001111111101010000); #20
	MCMC_indirect_write(11'd2030, 68'b11100110101110111101101001110010011100100110110010110101010010011101); #20
	MCMC_indirect_write(11'd2031, 68'b11111100011100000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2032, 68'b11011000100000011101111001111011001100010110111101111010111000100111); #20
	MCMC_indirect_write(11'd2033, 68'b10000000000000000111111101011000011111001100111001011101010010010010); #20
	MCMC_indirect_write(11'd2034, 68'b01111001100011111100111010101001101001000100001111110110001010110111); #20
	MCMC_indirect_write(11'd2035, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2036, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2037, 68'b11110011111010100111110010001000001101110100000001111100100001000101); #20
	MCMC_indirect_write(11'd2038, 68'b10000000000000000100000000000000001000000000000000011011000000111001); #20
	MCMC_indirect_write(11'd2039, 68'b11100010011101110110101101010000101101011111010111111001010010010111); #20
	MCMC_indirect_write(11'd2040, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2041, 68'b10000000000000000100000000000000001000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2042, 68'b10100100101011101110010111110001001101111110111100111101001000010011); #20
	MCMC_indirect_write(11'd2043, 68'b10111011110100110101010101101110111011111000000101110101011111111011); #20
	MCMC_indirect_write(11'd2044, 68'b11100011011011000110111000011001111000000000000000010000000000000000); #20
	MCMC_indirect_write(11'd2045, 68'b11010011101110001110000100011101111111010010001000011001001011101110); #20
	MCMC_indirect_write(11'd2046, 68'b10001111000011001100100001101001010111011011100001010000010111011001); #20
	MCMC_indirect_write(11'd2047, 68'b10111001111011111100110111000110101000101100101111110100010010000010); #20

	//start core (address = 5 in define)
	apb_write(`START_ADDR, 1);
	


	#10000 $finish;
	
	//	Test for 256 signals
	//	FIFO_indirect_write(8'b00000000, 18'b110001000010000001); #20
	//	FIFO_indirect_write(8'b00000001, 18'b001000100000100101); #20
	//	FIFO_indirect_write(8'b00000010, 18'b000011100110101111); #20
	//	FIFO_indirect_write(8'b00000011, 18'b101001110010100000); #20
	//	FIFO_indirect_write(8'd4, 18'b001001000101010101); #20
	//	FIFO_indirect_write(8'd5, 18'b001001100000010011); #20
	//	FIFO_indirect_write(8'd6, 18'b101011111111011110); #20
	//	FIFO_indirect_write(8'd7, 18'b100001001000101000); #20
	//	FIFO_indirect_write(8'd8, 18'b110100110010100011); #20
	//	FIFO_indirect_write(8'd9, 18'b100100101001110001); #20
	//	FIFO_indirect_write(8'd10, 18'b101100011000100111); #20
	//	FIFO_indirect_write(8'd11, 18'b000010011111001010); #20
	//	FIFO_indirect_write(8'd12, 18'b111110110110101100); #20
	//	FIFO_indirect_write(8'd13, 18'b011101000011001110); #20
	//	FIFO_indirect_write(8'd14, 18'b001100011100110101); #20
	//	FIFO_indirect_write(8'd15, 18'b011100111010011001); #20
	//	FIFO_indirect_write(8'd16, 18'b011000001010111010); #20
	//	FIFO_indirect_write(8'd17, 18'b111111010111010010); #20
	//	FIFO_indirect_write(8'd18, 18'b011010001100001011); #20
	//	FIFO_indirect_write(8'd19, 18'b000110010100011110); #20
	//	FIFO_indirect_write(8'd20, 18'b001100010101111111); #20
	//	FIFO_indirect_write(8'd21, 18'b111111000010001011); #20
	//	FIFO_indirect_write(8'd22, 18'b010011010000011000); #20
	//	FIFO_indirect_write(8'd23, 18'b000101000100010101); #20
	//	FIFO_indirect_write(8'd24, 18'b101001110110011010); #20
	//	FIFO_indirect_write(8'd25, 18'b101010100001010011); #20
	//	FIFO_indirect_write(8'd26, 18'b111101101010000111); #20
	//	FIFO_indirect_write(8'd27, 18'b001100111110100101); #20
	//	FIFO_indirect_write(8'd28, 18'b110101111000000110); #20
	//	FIFO_indirect_write(8'd29, 18'b111100011011110000); #20
	//	FIFO_indirect_write(8'd30, 18'b001010001000000000); #20
	//	FIFO_indirect_write(8'd31, 18'b101001000110001110); #20
	//	FIFO_indirect_write(8'd32, 18'b111111110000000001); #20
	//	FIFO_indirect_write(8'd33, 18'b010000000010010100); #20
	//	FIFO_indirect_write(8'd34, 18'b011001000101100100); #20
	//	FIFO_indirect_write(8'd35, 18'b010110100110111110); #20
	//	FIFO_indirect_write(8'd36, 18'b001100101110100111); #20
	//	FIFO_indirect_write(8'd37, 18'b001011100111000010); #20
	//	FIFO_indirect_write(8'd38, 18'b000000010101001011); #20
	//	FIFO_indirect_write(8'd39, 18'b100001100111101100); #20
	//	FIFO_indirect_write(8'd40, 18'b010110001001000101); #20
	//	FIFO_indirect_write(8'd41, 18'b100111001001011111); #20
	//	FIFO_indirect_write(8'd42, 18'b010101111000010000); #20
	//	FIFO_indirect_write(8'd43, 18'b101011010111101101); #20
	//	FIFO_indirect_write(8'd44, 18'b001101101111011000); #20
	//	FIFO_indirect_write(8'd45, 18'b001001000011101010); #20
	//	FIFO_indirect_write(8'd46, 18'b000011100110000000); #20
	//	FIFO_indirect_write(8'd47, 18'b000000101101100101); #20
	//	FIFO_indirect_write(8'd48, 18'b010111111010100100); #20
	//	FIFO_indirect_write(8'd49, 18'b111010100011001001); #20
	//	FIFO_indirect_write(8'd50, 18'b000010011101001110); #20
	//	FIFO_indirect_write(8'd51, 18'b000101001011101110); #20
	//	FIFO_indirect_write(8'd52, 18'b000101011110101010); #20
	//	FIFO_indirect_write(8'd53, 18'b011101111101101000); #20
	//	FIFO_indirect_write(8'd54, 18'b110111000101011011); #20
	//	FIFO_indirect_write(8'd55, 18'b011100110000101010); #20
	//	FIFO_indirect_write(8'd56, 18'b000110001100111011); #20
	//	FIFO_indirect_write(8'd57, 18'b010111011100101010); #20
	//	FIFO_indirect_write(8'd58, 18'b101001000101000110); #20
	//	FIFO_indirect_write(8'd59, 18'b110011011010111010); #20
	//	FIFO_indirect_write(8'd60, 18'b110001000011011100); #20
	//	FIFO_indirect_write(8'd61, 18'b111000010001100011); #20
	//	FIFO_indirect_write(8'd62, 18'b010111100111011001); #20
	//	FIFO_indirect_write(8'd63, 18'b110000111011100111); #20
	//	FIFO_indirect_write(8'd64, 18'b111101001001110101); #20
	//	FIFO_indirect_write(8'd65, 18'b011011110000001011); #20
	//	FIFO_indirect_write(8'd66, 18'b100010011101001010); #20
	//	FIFO_indirect_write(8'd67, 18'b101111010000000101); #20
	//	FIFO_indirect_write(8'd68, 18'b101110111001101011); #20
	//	FIFO_indirect_write(8'd69, 18'b101111100111001111); #20
	//	FIFO_indirect_write(8'd70, 18'b101111111011011100); #20
	//	FIFO_indirect_write(8'd71, 18'b001001001101101010); #20
	//	FIFO_indirect_write(8'd72, 18'b000101100001111010); #20
	//	FIFO_indirect_write(8'd73, 18'b000001100000000111); #20
	//	FIFO_indirect_write(8'd74, 18'b000110011101101001); #20
	//	FIFO_indirect_write(8'd75, 18'b010001111011100111); #20
	//	FIFO_indirect_write(8'd76, 18'b110001101110110111); #20
	//	FIFO_indirect_write(8'd77, 18'b011011100000111000); #20
	//	FIFO_indirect_write(8'd78, 18'b110001011000000000); #20
	//	FIFO_indirect_write(8'd79, 18'b100000100100100100); #20
	//	FIFO_indirect_write(8'd80, 18'b000100010100111001); #20
	//	FIFO_indirect_write(8'd81, 18'b101101001100010100); #20
	//	FIFO_indirect_write(8'd82, 18'b110110110011011111); #20
	//	FIFO_indirect_write(8'd83, 18'b011010111010011011); #20
	//	FIFO_indirect_write(8'd84, 18'b100001010111110011); #20
	//	FIFO_indirect_write(8'd85, 18'b110010111101101100); #20
	//	FIFO_indirect_write(8'd86, 18'b101110000110011101); #20
	//	FIFO_indirect_write(8'd87, 18'b010100011101011111); #20
	//	FIFO_indirect_write(8'd88, 18'b101100000110111111); #20
	//	FIFO_indirect_write(8'd89, 18'b011011011110110111); #20
	//	FIFO_indirect_write(8'd90, 18'b001101000011100101); #20
	//	FIFO_indirect_write(8'd91, 18'b101101110111001010); #20
	//	FIFO_indirect_write(8'd92, 18'b011001110011111000); #20
	//	FIFO_indirect_write(8'd93, 18'b010010110110001101); #20
	//	FIFO_indirect_write(8'd94, 18'b101011101000111111); #20
	//	FIFO_indirect_write(8'd95, 18'b111100010001000001); #20
	//	FIFO_indirect_write(8'd96, 18'b011101101001111111); #20
	//	FIFO_indirect_write(8'd97, 18'b110101011110000011); #20
	//	FIFO_indirect_write(8'd98, 18'b001001110001010011); #20
	//	FIFO_indirect_write(8'd99, 18'b101010000000000110); #20
	//	FIFO_indirect_write(8'd100, 18'b011101000101000010); #20
	//	FIFO_indirect_write(8'd101, 18'b101010110101001111); #20
	//	FIFO_indirect_write(8'd102, 18'b110110001110011001); #20
	//	FIFO_indirect_write(8'd103, 18'b110110011001101101); #20
	//	FIFO_indirect_write(8'd104, 18'b101001011101000000); #20
	//	FIFO_indirect_write(8'd105, 18'b110000111000010000); #20
	//	FIFO_indirect_write(8'd106, 18'b001000010010100100); #20
	//	FIFO_indirect_write(8'd107, 18'b001000001011000100); #20
	//	FIFO_indirect_write(8'd108, 18'b111000000100101111); #20
	//	FIFO_indirect_write(8'd109, 18'b011001011100010101); #20
	//	FIFO_indirect_write(8'd110, 18'b011110001101110110); #20
	//	FIFO_indirect_write(8'd111, 18'b101001011011101010); #20
	//	FIFO_indirect_write(8'd112, 18'b010010111110110011); #20
	//	FIFO_indirect_write(8'd113, 18'b011101010000101011); #20
	//	FIFO_indirect_write(8'd114, 18'b001100011111100111); #20
	//	FIFO_indirect_write(8'd115, 18'b100111101111110100); #20
	//	FIFO_indirect_write(8'd116, 18'b010110011111001100); #20
	//	FIFO_indirect_write(8'd117, 18'b110101001000110101); #20
	//	FIFO_indirect_write(8'd118, 18'b110100001001101101); #20
	//	FIFO_indirect_write(8'd119, 18'b011001000011010100); #20
	//	FIFO_indirect_write(8'd120, 18'b011000100001101010); #20
	//	FIFO_indirect_write(8'd121, 18'b010011001111010110); #20
	//	FIFO_indirect_write(8'd122, 18'b010000001000011111); #20
	//	FIFO_indirect_write(8'd123, 18'b110011010111101110); #20
	//	FIFO_indirect_write(8'd124, 18'b000001011011011111); #20
	//	FIFO_indirect_write(8'd125, 18'b001000010001101000); #20
	//	FIFO_indirect_write(8'd126, 18'b110111011000110100); #20
	//	FIFO_indirect_write(8'd127, 18'b000001100111100101); #20
	//	FIFO_indirect_write(8'd128, 18'b010110001101100110); #20
	//	FIFO_indirect_write(8'd129, 18'b111101110111110111); #20
	//	FIFO_indirect_write(8'd130, 18'b010100000001101010); #20
	//	FIFO_indirect_write(8'd131, 18'b111000110110111100); #20
	//	FIFO_indirect_write(8'd132, 18'b001011000011011010); #20
	//	FIFO_indirect_write(8'd133, 18'b111000011001011101); #20
	//	FIFO_indirect_write(8'd134, 18'b110101010110011110); #20
	//	FIFO_indirect_write(8'd135, 18'b001100111010110010); #20
	//	FIFO_indirect_write(8'd136, 18'b010100010111001111); #20
	//	FIFO_indirect_write(8'd137, 18'b000100101110000110); #20
	//	FIFO_indirect_write(8'd138, 18'b011101100100001000); #20
	//	FIFO_indirect_write(8'd139, 18'b101111011101001110); #20
	//	FIFO_indirect_write(8'd140, 18'b100010110011100000); #20
	//	FIFO_indirect_write(8'd141, 18'b011000111010001011); #20
	//	FIFO_indirect_write(8'd142, 18'b101001010011011100); #20
	//	FIFO_indirect_write(8'd143, 18'b011010100001011010); #20
	//	FIFO_indirect_write(8'd144, 18'b010101110100110101); #20
	//	FIFO_indirect_write(8'd145, 18'b110100011111001100); #20
	//	FIFO_indirect_write(8'd146, 18'b010010100001101111); #20
	//	FIFO_indirect_write(8'd147, 18'b100010011010000011); #20
	//	FIFO_indirect_write(8'd148, 18'b011000001110011110); #20
	//	FIFO_indirect_write(8'd149, 18'b101001011000010000); #20
	//	FIFO_indirect_write(8'd150, 18'b001011110010110101); #20
	//	FIFO_indirect_write(8'd151, 18'b110110010000010111); #20
	//	FIFO_indirect_write(8'd152, 18'b000000001001101100); #20
	//	FIFO_indirect_write(8'd153, 18'b100101111000011001); #20
	//	FIFO_indirect_write(8'd154, 18'b111011000100010010); #20
	//	FIFO_indirect_write(8'd155, 18'b010000110101110010); #20
	//	FIFO_indirect_write(8'd156, 18'b011110011000001010); #20
	//	FIFO_indirect_write(8'd157, 18'b000100001111111011); #20
	//	FIFO_indirect_write(8'd158, 18'b101110110000100011); #20
	//	FIFO_indirect_write(8'd159, 18'b011111010000100011); #20
	//	FIFO_indirect_write(8'd160, 18'b010001011011100001); #20
	//	FIFO_indirect_write(8'd161, 18'b000000010011011100); #20
	//	FIFO_indirect_write(8'd162, 18'b110101111110011010); #20
	//	FIFO_indirect_write(8'd163, 18'b101110111001010111); #20
	//	FIFO_indirect_write(8'd164, 18'b011001001111111101); #20
	//	FIFO_indirect_write(8'd165, 18'b111101001101101010); #20
	//	FIFO_indirect_write(8'd166, 18'b110111000100110110); #20
	//	FIFO_indirect_write(8'd167, 18'b110010101010000101); #20
	//	FIFO_indirect_write(8'd168, 18'b001101100111110000); #20
	//	FIFO_indirect_write(8'd169, 18'b010000100011111111); #20
	//	FIFO_indirect_write(8'd170, 18'b100100101010110110); #20
	//	FIFO_indirect_write(8'd171, 18'b011101100111001010); #20
	//	FIFO_indirect_write(8'd172, 18'b011000100101101110); #20
	//	FIFO_indirect_write(8'd173, 18'b100000100011010110); #20
	//	FIFO_indirect_write(8'd174, 18'b001010101110010000); #20
	//	FIFO_indirect_write(8'd175, 18'b001100100101100010); #20
	//	FIFO_indirect_write(8'd176, 18'b001101001100000001); #20
	//	FIFO_indirect_write(8'd177, 18'b000110100101011110); #20
	//	FIFO_indirect_write(8'd178, 18'b100000110100011111); #20
	//	FIFO_indirect_write(8'd179, 18'b111010001000001110); #20
	//	FIFO_indirect_write(8'd180, 18'b110010000100010000); #20
	//	FIFO_indirect_write(8'd181, 18'b011001110000101101); #20
	//	FIFO_indirect_write(8'd182, 18'b010111100101110001); #20
	//	FIFO_indirect_write(8'd183, 18'b010011000001110000); #20
	//	FIFO_indirect_write(8'd184, 18'b110110000110110011); #20
	//	FIFO_indirect_write(8'd185, 18'b110111110101101111); #20
	//	FIFO_indirect_write(8'd186, 18'b000101101010011110); #20
	//	FIFO_indirect_write(8'd187, 18'b010011000100010010); #20
	//	FIFO_indirect_write(8'd188, 18'b000111100110010010); #20
	//	FIFO_indirect_write(8'd189, 18'b011111010001110111); #20
	//	FIFO_indirect_write(8'd190, 18'b011110100001110101); #20
	//	FIFO_indirect_write(8'd191, 18'b011001100100111100); #20
	//	FIFO_indirect_write(8'd192, 18'b110011010100001101); #20
	//	FIFO_indirect_write(8'd193, 18'b100011001110111001); #20
	//	FIFO_indirect_write(8'd194, 18'b011011001000000110); #20
	//	FIFO_indirect_write(8'd195, 18'b111110100100111101); #20
	//	FIFO_indirect_write(8'd196, 18'b110000000010010110); #20
	//	FIFO_indirect_write(8'd197, 18'b101111011001110111); #20
	//	FIFO_indirect_write(8'd198, 18'b111101010000100010); #20
	//	FIFO_indirect_write(8'd199, 18'b011011010001111001); #20
	//	FIFO_indirect_write(8'd200, 18'b001000011101101001); #20
	//	FIFO_indirect_write(8'd201, 18'b000101100111010011); #20
	//	FIFO_indirect_write(8'd202, 18'b011111010001001110); #20
	//	FIFO_indirect_write(8'd203, 18'b000000010101000011); #20
	//	FIFO_indirect_write(8'd204, 18'b000001011110001001); #20
	//	FIFO_indirect_write(8'd205, 18'b111001000000011001); #20
	//	FIFO_indirect_write(8'd206, 18'b010110001010010000); #20
	//	FIFO_indirect_write(8'd207, 18'b101110000010100001); #20
	//	FIFO_indirect_write(8'd208, 18'b100000010111000100); #20
	//	FIFO_indirect_write(8'd209, 18'b110010001111001110); #20
	//	FIFO_indirect_write(8'd210, 18'b011110101000111100); #20
	//	FIFO_indirect_write(8'd211, 18'b101111011000100110); #20
	//	FIFO_indirect_write(8'd212, 18'b001111110011010111); #20
	//	FIFO_indirect_write(8'd213, 18'b011110011111001111); #20
	//	FIFO_indirect_write(8'd214, 18'b110110101000010010); #20
	//	FIFO_indirect_write(8'd215, 18'b000110101110101111); #20
	//	FIFO_indirect_write(8'd216, 18'b111010101111110101); #20
	//	FIFO_indirect_write(8'd217, 18'b111100010111100000); #20
	//	FIFO_indirect_write(8'd218, 18'b101100111001100000); #20
	//	FIFO_indirect_write(8'd219, 18'b110111000100010001); #20
	//	FIFO_indirect_write(8'd220, 18'b000111100000110111); #20
	//	FIFO_indirect_write(8'd221, 18'b111011111010100010); #20
	//	FIFO_indirect_write(8'd222, 18'b001110001010000111); #20
	//	FIFO_indirect_write(8'd223, 18'b111110010100011100); #20
	//	FIFO_indirect_write(8'd224, 18'b011010001111010010); #20
	//	FIFO_indirect_write(8'd225, 18'b101010010100011111); #20
	//	FIFO_indirect_write(8'd226, 18'b000011010101101001); #20
	//	FIFO_indirect_write(8'd227, 18'b111101000010010011); #20
	//	FIFO_indirect_write(8'd228, 18'b010000100101001111); #20
	//	FIFO_indirect_write(8'd229, 18'b100001110111010010); #20
	//	FIFO_indirect_write(8'd230, 18'b000110100110001000); #20
	//	FIFO_indirect_write(8'd231, 18'b110100111001111101); #20
	//	FIFO_indirect_write(8'd232, 18'b011111101000000010); #20
	//	FIFO_indirect_write(8'd233, 18'b111101111001111000); #20
	//	FIFO_indirect_write(8'd234, 18'b101000001000111011); #20
	//	FIFO_indirect_write(8'd235, 18'b100010101000100010); #20
	//	FIFO_indirect_write(8'd236, 18'b011011011101110001); #20
	//	FIFO_indirect_write(8'd237, 18'b100001000101110001); #20
	//	FIFO_indirect_write(8'd238, 18'b000100100001110010); #20
	//	FIFO_indirect_write(8'd239, 18'b110100000010010100); #20
	//	FIFO_indirect_write(8'd240, 18'b000001101111001001); #20
	//	FIFO_indirect_write(8'd241, 18'b010011100010001011); #20
	//	FIFO_indirect_write(8'd242, 18'b011010100101110001); #20
	//	FIFO_indirect_write(8'd243, 18'b000000101010011011); #20
	//	FIFO_indirect_write(8'd244, 18'b001011111110100110); #20
	//	FIFO_indirect_write(8'd245, 18'b011011011010000100); #20
	//	FIFO_indirect_write(8'd246, 18'b000000010001010001); #20
	//	FIFO_indirect_write(8'd247, 18'b100110101011101010); #20
	//	FIFO_indirect_write(8'd248, 18'b111010110110000001); #20
	//	FIFO_indirect_write(8'd249, 18'b011110000011100100); #20
	//	FIFO_indirect_write(8'd250, 18'b000011000101000110); #20
	//	FIFO_indirect_write(8'd251, 18'b000111110000011000); #20
	//	FIFO_indirect_write(8'd252, 18'b001000010100000111); #20
	//	FIFO_indirect_write(8'd253, 18'b100011000000001010); #20
	//	FIFO_indirect_write(8'd254, 18'b111000010000011001); #20
	//	FIFO_indirect_write(8'd255, 18'b010001111010011011); #20
	
	
	
end
endmodule